module SRAMTemplate(
  input         clock,
  input         reset,
  output        io_r_req_ready, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input         io_r_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [8:0]  io_r_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [28:0] io_r_resp_data_0_tag, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [1:0]  io_r_resp_data_0__type, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [38:0] io_r_resp_data_0_target, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output [2:0]  io_r_resp_data_0_brIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  output        io_r_resp_data_0_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input         io_w_req_valid, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [8:0]  io_w_req_bits_setIdx, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [28:0] io_w_req_bits_data_tag, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [1:0]  io_w_req_bits_data__type, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [38:0] io_w_req_bits_data_target, // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
  input  [2:0]  io_w_req_bits_data_brIdx // @[src/main/scala/utils/SRAMTemplate.scala 70:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [95:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [95:0] _RAND_10;
  reg [95:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] array_0_R0_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_R0_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_R0_clk; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [73:0] array_0_R0_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [8:0] array_0_W0_addr; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_W0_en; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire  array_0_W0_clk; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  wire [73:0] array_0_W0_data; // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
  reg  resetState; // @[src/main/scala/utils/SRAMTemplate.scala 80:30]
  reg [8:0] resetSet; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  wrap_wrap = resetSet == 9'h1ff; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [8:0] _wrap_value_T_1 = resetSet + 9'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  resetFinish = resetState & wrap_wrap; // @[src/main/scala/chisel3/util/Counter.scala 118:{16,23} 117:24]
  wire  _GEN_2 = resetFinish ? 1'h0 : resetState; // @[src/main/scala/utils/SRAMTemplate.scala 82:24 80:30 82:38]
  wire  wen = io_w_req_valid | resetState; // @[src/main/scala/utils/SRAMTemplate.scala 88:52]
  wire  _realRen_T = ~wen; // @[src/main/scala/utils/SRAMTemplate.scala 89:41]
  wire [73:0] _wdataword_T = {io_w_req_bits_data_tag,io_w_req_bits_data__type,io_w_req_bits_data_target,
    io_w_req_bits_data_brIdx,1'h1}; // @[src/main/scala/utils/SRAMTemplate.scala 92:78]
  reg  rdata_REG; // @[src/main/scala/utils/Hold.scala 28:106]
  reg [73:0] rdata_r_0; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [73:0] _GEN_14 = rdata_REG ? array_0_R0_data : rdata_r_0; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  resetState_p; // @[src/main/scala/utils/SRAMTemplate.scala 80:30]
  wire  resetState_t = resetState ^ resetState_p; // @[src/main/scala/utils/SRAMTemplate.scala 80:30]
  wire  toggle_0_clock;
  wire  toggle_0_reset;
  wire  toggle_0_valid;
  reg  toggle_0_valid_reg;
  reg [8:0] resetSet_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [8:0] resetSet_t = resetSet ^ resetSet_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  toggle_1_clock;
  wire  toggle_1_reset;
  wire [8:0] toggle_1_valid;
  reg [8:0] toggle_1_valid_reg;
  reg  rdata_REG_p; // @[src/main/scala/utils/Hold.scala 28:106]
  wire  rdata_REG_t = rdata_REG ^ rdata_REG_p; // @[src/main/scala/utils/Hold.scala 28:106]
  wire  toggle_10_clock;
  wire  toggle_10_reset;
  wire  toggle_10_valid;
  reg  toggle_10_valid_reg;
  reg [73:0] rdata_r_0_p; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [73:0] rdata_r_0_t = rdata_r_0 ^ rdata_r_0_p; // @[src/main/scala/utils/Hold.scala 23:65]
  wire  toggle_11_clock;
  wire  toggle_11_reset;
  wire [73:0] toggle_11_valid;
  reg [73:0] toggle_11_valid_reg;
  array_0 array_0 ( // @[src/main/scala/utils/SRAMTemplate.scala 76:26]
    .R0_addr(array_0_R0_addr),
    .R0_en(array_0_R0_en),
    .R0_clk(array_0_R0_clk),
    .R0_data(array_0_R0_data),
    .W0_addr(array_0_W0_addr),
    .W0_en(array_0_W0_en),
    .W0_clk(array_0_W0_clk),
    .W0_data(array_0_W0_data)
  );
  GEN_w1_toggle #(.COVER_INDEX(0)) toggle_0 (
    .clock(toggle_0_clock),
    .reset(toggle_0_reset),
    .valid(toggle_0_valid)
  );
  GEN_w9_toggle #(.COVER_INDEX(1)) toggle_1 (
    .clock(toggle_1_clock),
    .reset(toggle_1_reset),
    .valid(toggle_1_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10)) toggle_10 (
    .clock(toggle_10_clock),
    .reset(toggle_10_reset),
    .valid(toggle_10_valid)
  );
  GEN_w74_toggle #(.COVER_INDEX(11)) toggle_11 (
    .clock(toggle_11_clock),
    .reset(toggle_11_reset),
    .valid(toggle_11_valid)
  );
  assign io_r_req_ready = ~resetState & _realRen_T; // @[src/main/scala/utils/SRAMTemplate.scala 101:33]
  assign io_r_resp_data_0_tag = _GEN_14[73:45]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0__type = _GEN_14[44:43]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0_target = _GEN_14[42:4]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0_brIdx = _GEN_14[3:1]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign io_r_resp_data_0_valid = _GEN_14[0]; // @[src/main/scala/utils/SRAMTemplate.scala 98:78]
  assign array_0_R0_addr = io_r_req_bits_setIdx; // @[src/main/scala/utils/Hold.scala 28:87]
  assign array_0_R0_en = io_r_req_valid & ~wen; // @[src/main/scala/utils/SRAMTemplate.scala 89:38]
  assign array_0_R0_clk = clock; // @[src/main/scala/utils/Hold.scala 28:{87,87}]
  assign array_0_W0_addr = resetState ? resetSet : io_w_req_bits_setIdx; // @[src/main/scala/utils/SRAMTemplate.scala 91:19]
  assign array_0_W0_en = io_w_req_valid | resetState; // @[src/main/scala/utils/SRAMTemplate.scala 88:52]
  assign array_0_W0_clk = clock; // @[src/main/scala/utils/SRAMTemplate.scala 95:14]
  assign array_0_W0_data = resetState ? 74'h0 : _wdataword_T; // @[src/main/scala/utils/SRAMTemplate.scala 92:22]
  assign toggle_0_clock = clock;
  assign toggle_0_reset = reset;
  assign toggle_0_valid = resetState ^ toggle_0_valid_reg;
  assign toggle_1_clock = clock;
  assign toggle_1_reset = reset;
  assign toggle_1_valid = resetSet ^ toggle_1_valid_reg;
  assign toggle_10_clock = clock;
  assign toggle_10_reset = reset;
  assign toggle_10_valid = rdata_REG ^ toggle_10_valid_reg;
  assign toggle_11_clock = clock;
  assign toggle_11_reset = reset;
  assign toggle_11_valid = rdata_r_0 ^ toggle_11_valid_reg;
  always @(posedge clock) begin
    resetState <= reset | _GEN_2; // @[src/main/scala/utils/SRAMTemplate.scala 80:{30,30}]
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      resetSet <= 9'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (resetState) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      resetSet <= _wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    rdata_REG <= io_r_req_valid & ~wen; // @[src/main/scala/utils/SRAMTemplate.scala 89:38]
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      rdata_r_0 <= 74'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (rdata_REG) begin // @[src/main/scala/utils/Hold.scala 23:65]
      rdata_r_0 <= array_0_R0_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    resetState_p <= resetState; // @[src/main/scala/utils/SRAMTemplate.scala 80:30]
    toggle_0_valid_reg <= resetState;
    resetSet_p <= resetSet; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    toggle_1_valid_reg <= resetSet;
    rdata_REG_p <= rdata_REG; // @[src/main/scala/utils/Hold.scala 28:106]
    toggle_10_valid_reg <= rdata_REG;
    rdata_r_0_p <= rdata_r_0; // @[src/main/scala/utils/Hold.scala 23:65]
    toggle_11_valid_reg <= rdata_r_0;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  resetState = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  resetSet = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  rdata_REG = _RAND_2[0:0];
  _RAND_3 = {3{`RANDOM}};
  rdata_r_0 = _RAND_3[73:0];
  _RAND_4 = {1{`RANDOM}};
  resetState_p = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  toggle_0_valid_reg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  resetSet_p = _RAND_6[8:0];
  _RAND_7 = {1{`RANDOM}};
  toggle_1_valid_reg = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  rdata_REG_p = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  toggle_10_valid_reg = _RAND_9[0:0];
  _RAND_10 = {3{`RANDOM}};
  rdata_r_0_p = _RAND_10[73:0];
  _RAND_11 = {3{`RANDOM}};
  toggle_11_valid_reg = _RAND_11[73:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(resetState_t); // @[src/main/scala/utils/SRAMTemplate.scala 80:30]
    end
    //
    if (enToggle_past) begin
      cover(resetSet_t[0]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(resetSet_t[1]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(resetSet_t[2]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(resetSet_t[3]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(resetSet_t[4]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(resetSet_t[5]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(resetSet_t[6]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(resetSet_t[7]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(resetSet_t[8]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(rdata_REG_t); // @[src/main/scala/utils/Hold.scala 28:106]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[0]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[1]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[2]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[3]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[4]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[5]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[6]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[7]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[8]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[9]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[10]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[11]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[12]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[13]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[14]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[15]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[16]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[17]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[18]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[19]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[20]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[21]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[22]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[23]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[24]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[25]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[26]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[27]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[28]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[29]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[30]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[31]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[32]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[33]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[34]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[35]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[36]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[37]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[38]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[39]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[40]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[41]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[42]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[43]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[44]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[45]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[46]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[47]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[48]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[49]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[50]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[51]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[52]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[53]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[54]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[55]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[56]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[57]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[58]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[59]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[60]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[61]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[62]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[63]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[64]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[65]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[66]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[67]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[68]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[69]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[70]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[71]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[72]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[73]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
  end
endmodule
module BPU_inorder(
  input         clock,
  input         reset,
  input         io_in_pc_valid, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  input  [38:0] io_in_pc_bits, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  output [38:0] io_out_target, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  input         io_flush, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  output [2:0]  io_brIdx, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  output        io_crosslineJump, // @[src/main/scala/nutcore/frontend/BPU.scala 281:14]
  input         bpuUpdateReq_valid,
  input  [38:0] bpuUpdateReq_pc,
  input         bpuUpdateReq_isMissPredict,
  input  [38:0] bpuUpdateReq_actualTarget,
  input  [6:0]  bpuUpdateReq_fuOpType,
  input  [1:0]  bpuUpdateReq_btbType,
  input         bpuUpdateReq_isRVC,
  input         MOUFlushICache,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire  btb_clock; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_reset; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_io_r_req_ready; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_io_r_req_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [8:0] btb_io_r_req_bits_setIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [28:0] btb_io_r_resp_data_0_tag; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [1:0] btb_io_r_resp_data_0__type; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [38:0] btb_io_r_resp_data_0_target; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [2:0] btb_io_r_resp_data_0_brIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_io_r_resp_data_0_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire  btb_io_w_req_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [8:0] btb_io_w_req_bits_setIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [28:0] btb_io_w_req_bits_data_tag; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [1:0] btb_io_w_req_bits_data__type; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [38:0] btb_io_w_req_bits_data_target; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  wire [2:0] btb_io_w_req_bits_data_brIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
  reg [38:0] ras [0:15]; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire  ras_rasTarget_MPORT_en; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire [3:0] ras_rasTarget_MPORT_addr; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire [38:0] ras_rasTarget_MPORT_data; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire [38:0] ras_MPORT_1_data; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire [3:0] ras_MPORT_1_addr; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire  ras_MPORT_1_mask; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  wire  ras_MPORT_1_en; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  reg  flush; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = io_in_pc_valid ? 1'h0 : flush; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = io_flush | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [38:0] pcLatch; // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
  wire [28:0] btbRead_tag = btb_io_r_resp_data_0_tag; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire  btbRead_valid = btb_io_r_resp_data_0_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire  _btbHit_T_7 = btb_io_r_req_ready & btb_io_r_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  btbHit_REG; // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
  wire [2:0] btbRead_brIdx = btb_io_r_resp_data_0_brIdx; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire  btbHit = btbRead_valid & btbRead_tag == pcLatch[38:10] & ~flush & btbHit_REG & ~(pcLatch[1] & btbRead_brIdx[0]); // @[src/main/scala/nutcore/frontend/BPU.scala 320:131]
  wire  crosslineJump = btbRead_brIdx[2] & btbHit; // @[src/main/scala/nutcore/frontend/BPU.scala 327:40]
  wire [1:0] _T_9 = io_out_valid ? 2'h3 : 2'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 332:94]
  reg [3:0] sp_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [38:0] rasTarget; // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
  wire  _T_19 = ~bpuUpdateReq_pc[1]; // @[src/main/scala/nutcore/frontend/BPU.scala 353:150]
  wire  _btbWrite_brIdx_T_3 = bpuUpdateReq_pc[2:0] == 3'h6 & ~bpuUpdateReq_isRVC; // @[src/main/scala/nutcore/frontend/BPU.scala 367:46]
  wire [1:0] btbWrite_brIdx_hi = {_btbWrite_brIdx_T_3,bpuUpdateReq_pc[1]}; // @[src/main/scala/nutcore/frontend/BPU.scala 367:24]
  wire  _T_27 = bpuUpdateReq_fuOpType == 7'h5c; // @[src/main/scala/nutcore/frontend/BPU.scala 403:24]
  wire [3:0] _T_29 = sp_value + 4'h1; // @[src/main/scala/nutcore/frontend/BPU.scala 404:26]
  wire [38:0] _T_31 = bpuUpdateReq_pc + 39'h2; // @[src/main/scala/nutcore/frontend/BPU.scala 404:55]
  wire [38:0] _T_33 = bpuUpdateReq_pc + 39'h4; // @[src/main/scala/nutcore/frontend/BPU.scala 404:69]
  wire  _T_36 = sp_value == 4'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 409:21]
  wire [3:0] _value_T_4 = sp_value - 4'h1; // @[src/main/scala/nutcore/frontend/BPU.scala 412:53]
  wire [3:0] _value_T_5 = _T_36 ? 4'h0 : _value_T_4; // @[src/main/scala/nutcore/frontend/BPU.scala 412:22]
  wire [1:0] btbRead__type = btb_io_r_resp_data_0__type; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire [38:0] btbRead_target = btb_io_r_resp_data_0_target; // @[src/main/scala/nutcore/frontend/BPU.scala 315:21 316:11]
  wire [3:0] _io_brIdx_T_1 = {1'h1,crosslineJump,_T_9}; // @[src/main/scala/nutcore/frontend/BPU.scala 419:35]
  wire [3:0] _GEN_7 = {{1'd0}, btbRead_brIdx}; // @[src/main/scala/nutcore/frontend/BPU.scala 419:30]
  wire [3:0] _io_brIdx_T_2 = _GEN_7 & _io_brIdx_T_1; // @[src/main/scala/nutcore/frontend/BPU.scala 419:30]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  flush_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  flush_t = flush ^ flush_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_85_clock;
  wire  toggle_85_reset;
  wire  toggle_85_valid;
  reg  toggle_85_valid_reg;
  reg [38:0] pcLatch_p; // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
  wire [38:0] pcLatch_t = pcLatch ^ pcLatch_p; // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
  wire  toggle_86_clock;
  wire  toggle_86_reset;
  wire [38:0] toggle_86_valid;
  reg [38:0] toggle_86_valid_reg;
  reg  btbHit_REG_p; // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
  wire  btbHit_REG_t = btbHit_REG ^ btbHit_REG_p; // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
  wire  toggle_125_clock;
  wire  toggle_125_reset;
  wire  toggle_125_valid;
  reg  toggle_125_valid_reg;
  reg [3:0] sp_value_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [3:0] sp_value_t = sp_value ^ sp_value_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  toggle_126_clock;
  wire  toggle_126_reset;
  wire [3:0] toggle_126_valid;
  reg [3:0] toggle_126_valid_reg;
  reg [38:0] rasTarget_p; // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
  wire [38:0] rasTarget_t = rasTarget ^ rasTarget_p; // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
  wire  toggle_130_clock;
  wire  toggle_130_reset;
  wire [38:0] toggle_130_valid;
  reg [38:0] toggle_130_valid_reg;
  SRAMTemplate btb ( // @[src/main/scala/nutcore/frontend/BPU.scala 302:19]
    .clock(btb_clock),
    .reset(btb_reset),
    .io_r_req_ready(btb_io_r_req_ready),
    .io_r_req_valid(btb_io_r_req_valid),
    .io_r_req_bits_setIdx(btb_io_r_req_bits_setIdx),
    .io_r_resp_data_0_tag(btb_io_r_resp_data_0_tag),
    .io_r_resp_data_0__type(btb_io_r_resp_data_0__type),
    .io_r_resp_data_0_target(btb_io_r_resp_data_0_target),
    .io_r_resp_data_0_brIdx(btb_io_r_resp_data_0_brIdx),
    .io_r_resp_data_0_valid(btb_io_r_resp_data_0_valid),
    .io_w_req_valid(btb_io_w_req_valid),
    .io_w_req_bits_setIdx(btb_io_w_req_bits_setIdx),
    .io_w_req_bits_data_tag(btb_io_w_req_bits_data_tag),
    .io_w_req_bits_data__type(btb_io_w_req_bits_data__type),
    .io_w_req_bits_data_target(btb_io_w_req_bits_data_target),
    .io_w_req_bits_data_brIdx(btb_io_w_req_bits_data_brIdx)
  );
  GEN_w1_toggle #(.COVER_INDEX(85)) toggle_85 (
    .clock(toggle_85_clock),
    .reset(toggle_85_reset),
    .valid(toggle_85_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(86)) toggle_86 (
    .clock(toggle_86_clock),
    .reset(toggle_86_reset),
    .valid(toggle_86_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(125)) toggle_125 (
    .clock(toggle_125_clock),
    .reset(toggle_125_reset),
    .valid(toggle_125_valid)
  );
  GEN_w4_toggle #(.COVER_INDEX(126)) toggle_126 (
    .clock(toggle_126_clock),
    .reset(toggle_126_reset),
    .valid(toggle_126_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(130)) toggle_130 (
    .clock(toggle_130_clock),
    .reset(toggle_130_reset),
    .valid(toggle_130_valid)
  );
  assign ras_rasTarget_MPORT_en = 1'h1;
  assign ras_rasTarget_MPORT_addr = sp_value;
  assign ras_rasTarget_MPORT_data = ras[ras_rasTarget_MPORT_addr]; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
  assign ras_MPORT_1_data = bpuUpdateReq_isRVC ? _T_31 : _T_33;
  assign ras_MPORT_1_addr = sp_value + 4'h1;
  assign ras_MPORT_1_mask = 1'h1;
  assign ras_MPORT_1_en = bpuUpdateReq_valid & _T_27;
  assign io_out_target = btbRead__type == 2'h3 ? rasTarget : btbRead_target; // @[src/main/scala/nutcore/frontend/BPU.scala 416:23]
  assign io_out_valid = 1'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 420:16]
  assign io_brIdx = _io_brIdx_T_2[2:0]; // @[src/main/scala/nutcore/frontend/BPU.scala 419:13]
  assign io_crosslineJump = btbRead_brIdx[2] & btbHit; // @[src/main/scala/nutcore/frontend/BPU.scala 327:40]
  assign btb_clock = clock;
  assign btb_reset = reset | (MOUFlushICache | MOUFlushTLB); // @[src/main/scala/nutcore/frontend/BPU.scala 308:29]
  assign btb_io_r_req_valid = io_in_pc_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 311:22]
  assign btb_io_r_req_bits_setIdx = io_in_pc_bits[9:1]; // @[src/main/scala/nutcore/frontend/BPU.scala 35:65]
  assign btb_io_w_req_valid = bpuUpdateReq_isMissPredict & bpuUpdateReq_valid; // @[src/main/scala/nutcore/frontend/BPU.scala 375:43]
  assign btb_io_w_req_bits_setIdx = bpuUpdateReq_pc[9:1]; // @[src/main/scala/nutcore/frontend/BPU.scala 35:65]
  assign btb_io_w_req_bits_data_tag = bpuUpdateReq_pc[38:10]; // @[src/main/scala/nutcore/frontend/BPU.scala 35:65]
  assign btb_io_w_req_bits_data__type = bpuUpdateReq_btbType; // @[src/main/scala/nutcore/frontend/BPU.scala 349:21]
  assign btb_io_w_req_bits_data_target = bpuUpdateReq_actualTarget; // @[src/main/scala/nutcore/frontend/BPU.scala 349:21]
  assign btb_io_w_req_bits_data_brIdx = {btbWrite_brIdx_hi,_T_19}; // @[src/main/scala/nutcore/frontend/BPU.scala 367:24]
  assign toggle_85_clock = clock;
  assign toggle_85_reset = reset;
  assign toggle_85_valid = flush ^ toggle_85_valid_reg;
  assign toggle_86_clock = clock;
  assign toggle_86_reset = reset;
  assign toggle_86_valid = pcLatch ^ toggle_86_valid_reg;
  assign toggle_125_clock = clock;
  assign toggle_125_reset = reset;
  assign toggle_125_valid = btbHit_REG ^ toggle_125_valid_reg;
  assign toggle_126_clock = clock;
  assign toggle_126_reset = reset;
  assign toggle_126_valid = sp_value ^ toggle_126_valid_reg;
  assign toggle_130_clock = clock;
  assign toggle_130_reset = reset;
  assign toggle_130_valid = rasTarget ^ toggle_130_valid_reg;
  always @(posedge clock) begin
    if (ras_MPORT_1_en & ras_MPORT_1_mask) begin
      ras[ras_MPORT_1_addr] <= ras_MPORT_1_data; // @[src/main/scala/nutcore/frontend/BPU.scala 342:16]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      flush <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      flush <= _GEN_1;
    end
    if (io_in_pc_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
      pcLatch <= io_in_pc_bits; // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    if (reset) begin // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
      btbHit_REG <= 1'h0; // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
    end else begin
      btbHit_REG <= _btbHit_T_7; // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      sp_value <= 4'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (bpuUpdateReq_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 402:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[src/main/scala/nutcore/frontend/BPU.scala 403:45]
        sp_value <= _T_29; // @[src/main/scala/nutcore/frontend/BPU.scala 406:16]
      end else if (bpuUpdateReq_fuOpType == 7'h5e) begin // @[src/main/scala/nutcore/frontend/BPU.scala 408:48]
        sp_value <= _value_T_5; // @[src/main/scala/nutcore/frontend/BPU.scala 412:16]
      end
    end
    if (io_in_pc_valid) begin // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
      rasTarget <= ras_rasTarget_MPORT_data; // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    flush_p <= flush; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_85_valid_reg <= flush;
    pcLatch_p <= pcLatch; // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    toggle_86_valid_reg <= pcLatch;
    btbHit_REG_p <= btbHit_REG; // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
    toggle_125_valid_reg <= btbHit_REG;
    sp_value_p <= sp_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    toggle_126_valid_reg <= sp_value;
    rasTarget_p <= rasTarget; // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    toggle_130_valid_reg <= rasTarget;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ras[initvar] = _RAND_0[38:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  flush = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  pcLatch = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  btbHit_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  sp_value = _RAND_4[3:0];
  _RAND_5 = {2{`RANDOM}};
  rasTarget = _RAND_5[38:0];
  _RAND_6 = {1{`RANDOM}};
  flush_p = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  toggle_85_valid_reg = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  pcLatch_p = _RAND_8[38:0];
  _RAND_9 = {2{`RANDOM}};
  toggle_86_valid_reg = _RAND_9[38:0];
  _RAND_10 = {1{`RANDOM}};
  btbHit_REG_p = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  toggle_125_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  sp_value_p = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  toggle_126_valid_reg = _RAND_13[3:0];
  _RAND_14 = {2{`RANDOM}};
  rasTarget_p = _RAND_14[38:0];
  _RAND_15 = {2{`RANDOM}};
  toggle_130_valid_reg = _RAND_15[38:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(flush_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[0]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[1]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[2]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[3]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[4]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[5]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[6]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[7]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[8]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[9]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[10]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[11]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[12]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[13]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[14]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[15]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[16]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[17]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[18]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[19]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[20]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[21]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[22]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[23]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[24]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[25]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[26]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[27]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[28]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[29]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[30]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[31]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[32]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[33]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[34]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[35]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[36]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[37]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(pcLatch_t[38]); // @[src/main/scala/nutcore/frontend/BPU.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(btbHit_REG_t); // @[src/main/scala/nutcore/frontend/BPU.scala 320:93]
    end
    //
    if (enToggle_past) begin
      cover(sp_value_t[0]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(sp_value_t[1]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(sp_value_t[2]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(sp_value_t[3]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[0]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[1]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[2]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[3]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[4]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[5]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[6]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[7]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[8]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[9]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[10]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[11]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[12]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[13]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[14]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[15]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[16]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[17]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[18]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[19]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[20]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[21]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[22]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[23]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[24]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[25]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[26]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[27]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[28]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[29]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[30]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[31]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[32]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[33]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[34]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[35]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[36]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[37]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
    //
    if (enToggle_past) begin
      cover(rasTarget_t[38]); // @[src/main/scala/nutcore/frontend/BPU.scala 345:28]
    end
  end
endmodule
module IFU_inorder(
  input         clock,
  input         reset,
  input         io_imem_req_ready, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output        io_imem_req_valid, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [38:0] io_imem_req_bits_addr, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [81:0] io_imem_req_bits_user, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output        io_imem_resp_ready, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input         io_imem_resp_valid, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input  [63:0] io_imem_resp_bits_rdata, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input  [81:0] io_imem_resp_bits_user, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input         io_out_ready, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [63:0] io_out_bits_instr, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [38:0] io_out_bits_pc, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [38:0] io_out_bits_pnpc, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output        io_out_bits_exceptionVec_1, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [3:0]  io_out_bits_brIdx, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input  [38:0] io_redirect_target, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input         io_redirect_valid, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  output [3:0]  io_flushVec, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input         io_iaf, // @[src/main/scala/nutcore/frontend/IFU.scala 310:14]
  input         REG_valid,
  input  [38:0] REG_pc,
  input         REG_isMissPredict,
  input  [38:0] REG_actualTarget,
  input  [6:0]  REG_fuOpType,
  input  [1:0]  REG_btbType,
  input         REG_isRVC,
  input         flushICache,
  input         flushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  bp1_clock; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_reset; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_io_in_pc_valid; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [38:0] bp1_io_in_pc_bits; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [38:0] bp1_io_out_target; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_io_out_valid; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_io_flush; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [2:0] bp1_io_brIdx; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_io_crosslineJump; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_bpuUpdateReq_valid; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [38:0] bp1_bpuUpdateReq_pc; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_bpuUpdateReq_isMissPredict; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [38:0] bp1_bpuUpdateReq_actualTarget; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [6:0] bp1_bpuUpdateReq_fuOpType; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire [1:0] bp1_bpuUpdateReq_btbType; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_bpuUpdateReq_isRVC; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_MOUFlushICache; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  wire  bp1_MOUFlushTLB; // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
  reg [38:0] pc; // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
  wire  _pcUpdate_T = io_imem_req_ready & io_imem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  pcUpdate = io_redirect_valid | _pcUpdate_T; // @[src/main/scala/nutcore/frontend/IFU.scala 324:36]
  wire [38:0] _snpc_T_2 = pc + 39'h2; // @[src/main/scala/nutcore/frontend/IFU.scala 325:28]
  wire [38:0] _snpc_T_4 = pc + 39'h4; // @[src/main/scala/nutcore/frontend/IFU.scala 325:38]
  wire [38:0] snpc = pc[1] ? _snpc_T_2 : _snpc_T_4; // @[src/main/scala/nutcore/frontend/IFU.scala 325:17]
  reg  crosslineJumpLatch; // @[src/main/scala/nutcore/frontend/IFU.scala 330:35]
  reg [38:0] crosslineJumpTarget; // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
  wire [38:0] _npc_T_1 = crosslineJumpLatch ? crosslineJumpTarget : snpc; // @[src/main/scala/nutcore/frontend/IFU.scala 341:59]
  wire [38:0] npc = io_redirect_valid ? io_redirect_target : _npc_T_1; // @[src/main/scala/nutcore/frontend/IFU.scala 341:16]
  wire  _npcIsSeq_T_2 = crosslineJumpLatch ? 1'h0 : 1'h1; // @[src/main/scala/nutcore/frontend/IFU.scala 342:54]
  wire  npcIsSeq = io_redirect_valid ? 1'h0 : _npcIsSeq_T_2; // @[src/main/scala/nutcore/frontend/IFU.scala 342:21]
  wire [2:0] _brIdx_T = io_redirect_valid ? 3'h0 : bp1_io_brIdx; // @[src/main/scala/nutcore/frontend/IFU.scala 350:29]
  wire [42:0] x8_hi = {npcIsSeq,_brIdx_T,npc}; // @[src/main/scala/nutcore/frontend/IFU.scala 372:82]
  wire  _T_3 = io_imem_resp_ready & io_imem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_3 = io_imem_req_valid | r; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _T_4 = |io_flushVec; // @[src/main/scala/nutcore/frontend/IFU.scala 396:37]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [38:0] pc_p; // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
  wire [38:0] pc_t = pc ^ pc_p; // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
  wire  toggle_169_clock;
  wire  toggle_169_reset;
  wire [38:0] toggle_169_valid;
  reg [38:0] toggle_169_valid_reg;
  reg  crosslineJumpLatch_p; // @[src/main/scala/nutcore/frontend/IFU.scala 330:35]
  wire  crosslineJumpLatch_t = crosslineJumpLatch ^ crosslineJumpLatch_p; // @[src/main/scala/nutcore/frontend/IFU.scala 330:35]
  wire  toggle_208_clock;
  wire  toggle_208_reset;
  wire  toggle_208_valid;
  reg  toggle_208_valid_reg;
  reg [38:0] crosslineJumpTarget_p; // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
  wire [38:0] crosslineJumpTarget_t = crosslineJumpTarget ^ crosslineJumpTarget_p; // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
  wire  toggle_209_clock;
  wire  toggle_209_reset;
  wire [38:0] toggle_209_valid;
  reg [38:0] toggle_209_valid_reg;
  reg  r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  r_t = r ^ r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_248_clock;
  wire  toggle_248_reset;
  wire  toggle_248_valid;
  reg  toggle_248_valid_reg;
  BPU_inorder bp1 ( // @[src/main/scala/nutcore/frontend/IFU.scala 327:19]
    .clock(bp1_clock),
    .reset(bp1_reset),
    .io_in_pc_valid(bp1_io_in_pc_valid),
    .io_in_pc_bits(bp1_io_in_pc_bits),
    .io_out_target(bp1_io_out_target),
    .io_out_valid(bp1_io_out_valid),
    .io_flush(bp1_io_flush),
    .io_brIdx(bp1_io_brIdx),
    .io_crosslineJump(bp1_io_crosslineJump),
    .bpuUpdateReq_valid(bp1_bpuUpdateReq_valid),
    .bpuUpdateReq_pc(bp1_bpuUpdateReq_pc),
    .bpuUpdateReq_isMissPredict(bp1_bpuUpdateReq_isMissPredict),
    .bpuUpdateReq_actualTarget(bp1_bpuUpdateReq_actualTarget),
    .bpuUpdateReq_fuOpType(bp1_bpuUpdateReq_fuOpType),
    .bpuUpdateReq_btbType(bp1_bpuUpdateReq_btbType),
    .bpuUpdateReq_isRVC(bp1_bpuUpdateReq_isRVC),
    .MOUFlushICache(bp1_MOUFlushICache),
    .MOUFlushTLB(bp1_MOUFlushTLB)
  );
  GEN_w39_toggle #(.COVER_INDEX(169)) toggle_169 (
    .clock(toggle_169_clock),
    .reset(toggle_169_reset),
    .valid(toggle_169_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(208)) toggle_208 (
    .clock(toggle_208_clock),
    .reset(toggle_208_reset),
    .valid(toggle_208_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(209)) toggle_209 (
    .clock(toggle_209_clock),
    .reset(toggle_209_reset),
    .valid(toggle_209_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(248)) toggle_248 (
    .clock(toggle_248_clock),
    .reset(toggle_248_reset),
    .valid(toggle_248_valid)
  );
  assign io_imem_req_valid = io_out_ready; // @[src/main/scala/nutcore/frontend/IFU.scala 373:21]
  assign io_imem_req_bits_addr = {pc[38:1],1'h0}; // @[src/main/scala/nutcore/frontend/IFU.scala 371:36]
  assign io_imem_req_bits_user = {x8_hi,pc}; // @[src/main/scala/nutcore/frontend/IFU.scala 372:82]
  assign io_imem_resp_ready = io_out_ready | io_flushVec[0]; // @[src/main/scala/nutcore/frontend/IFU.scala 375:38]
  assign io_out_valid = io_imem_resp_valid & ~io_flushVec[0]; // @[src/main/scala/nutcore/frontend/IFU.scala 393:38]
  assign io_out_bits_instr = io_imem_resp_bits_rdata; // @[src/main/scala/nutcore/frontend/IFU.scala 385:21]
  assign io_out_bits_pc = io_imem_resp_bits_user[38:0]; // @[src/main/scala/nutcore/frontend/IFU.scala 387:24]
  assign io_out_bits_pnpc = io_imem_resp_bits_user[77:39]; // @[src/main/scala/nutcore/frontend/IFU.scala 388:26]
  assign io_out_bits_exceptionVec_1 = io_iaf; // @[src/main/scala/nutcore/frontend/IFU.scala 392:46]
  assign io_out_bits_brIdx = io_imem_resp_bits_user[81:78]; // @[src/main/scala/nutcore/frontend/IFU.scala 389:27]
  assign io_flushVec = io_redirect_valid ? 4'hf : 4'h0; // @[src/main/scala/nutcore/frontend/IFU.scala 368:21]
  assign bp1_clock = clock;
  assign bp1_reset = reset;
  assign bp1_io_in_pc_valid = io_imem_req_ready & io_imem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  assign bp1_io_in_pc_bits = io_redirect_valid ? io_redirect_target : _npc_T_1; // @[src/main/scala/nutcore/frontend/IFU.scala 341:16]
  assign bp1_io_flush = io_redirect_valid; // @[src/main/scala/nutcore/frontend/IFU.scala 359:16]
  assign bp1_bpuUpdateReq_valid = REG_valid;
  assign bp1_bpuUpdateReq_pc = REG_pc;
  assign bp1_bpuUpdateReq_isMissPredict = REG_isMissPredict;
  assign bp1_bpuUpdateReq_actualTarget = REG_actualTarget;
  assign bp1_bpuUpdateReq_fuOpType = REG_fuOpType;
  assign bp1_bpuUpdateReq_btbType = REG_btbType;
  assign bp1_bpuUpdateReq_isRVC = REG_isRVC;
  assign bp1_MOUFlushICache = flushICache;
  assign bp1_MOUFlushTLB = flushTLB;
  assign toggle_169_clock = clock;
  assign toggle_169_reset = reset;
  assign toggle_169_valid = pc ^ toggle_169_valid_reg;
  assign toggle_208_clock = clock;
  assign toggle_208_reset = reset;
  assign toggle_208_valid = crosslineJumpLatch ^ toggle_208_valid_reg;
  assign toggle_209_clock = clock;
  assign toggle_209_reset = reset;
  assign toggle_209_valid = crosslineJumpTarget ^ toggle_209_valid_reg;
  assign toggle_248_clock = clock;
  assign toggle_248_reset = reset;
  assign toggle_248_valid = r ^ toggle_248_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
      pc <= 39'h80000000; // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end else if (pcUpdate) begin // @[src/main/scala/nutcore/frontend/IFU.scala 361:19]
      if (io_redirect_valid) begin // @[src/main/scala/nutcore/frontend/IFU.scala 341:16]
        pc <= io_redirect_target;
      end else if (crosslineJumpLatch) begin // @[src/main/scala/nutcore/frontend/IFU.scala 341:59]
        pc <= crosslineJumpTarget;
      end else begin
        pc <= snpc;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/frontend/IFU.scala 330:35]
      crosslineJumpLatch <= 1'h0; // @[src/main/scala/nutcore/frontend/IFU.scala 330:35]
    end else if (pcUpdate | bp1_io_flush) begin // @[src/main/scala/nutcore/frontend/IFU.scala 331:34]
      if (bp1_io_flush) begin // @[src/main/scala/nutcore/frontend/IFU.scala 332:30]
        crosslineJumpLatch <= 1'h0;
      end else begin
        crosslineJumpLatch <= bp1_io_crosslineJump & ~crosslineJumpLatch;
      end
    end
    if (bp1_io_crosslineJump) begin // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
      crosslineJumpTarget <= bp1_io_out_target; // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (_T_3) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      r <= _GEN_3;
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    pc_p <= pc; // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    toggle_169_valid_reg <= pc;
    crosslineJumpLatch_p <= crosslineJumpLatch; // @[src/main/scala/nutcore/frontend/IFU.scala 330:35]
    toggle_208_valid_reg <= crosslineJumpLatch;
    crosslineJumpTarget_p <= crosslineJumpTarget; // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    toggle_209_valid_reg <= crosslineJumpTarget;
    r_p <= r; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_248_valid_reg <= r;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc = _RAND_0[38:0];
  _RAND_1 = {1{`RANDOM}};
  crosslineJumpLatch = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  crosslineJumpTarget = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  r = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  pc_p = _RAND_4[38:0];
  _RAND_5 = {2{`RANDOM}};
  toggle_169_valid_reg = _RAND_5[38:0];
  _RAND_6 = {1{`RANDOM}};
  crosslineJumpLatch_p = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  toggle_208_valid_reg = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  crosslineJumpTarget_p = _RAND_8[38:0];
  _RAND_9 = {2{`RANDOM}};
  toggle_209_valid_reg = _RAND_9[38:0];
  _RAND_10 = {1{`RANDOM}};
  r_p = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  toggle_248_valid_reg = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(pc_t[0]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[1]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[2]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[3]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[4]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[5]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[6]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[7]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[8]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[9]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[10]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[11]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[12]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[13]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[14]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[15]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[16]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[17]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[18]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[19]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[20]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[21]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[22]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[23]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[24]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[25]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[26]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[27]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[28]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[29]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[30]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[31]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[32]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[33]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[34]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[35]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[36]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[37]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(pc_t[38]); // @[src/main/scala/nutcore/frontend/IFU.scala 323:19]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpLatch_t); // @[src/main/scala/nutcore/frontend/IFU.scala 330:35]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[0]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[1]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[2]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[3]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[4]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[5]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[6]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[7]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[8]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[9]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[10]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[11]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[12]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[13]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[14]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[15]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[16]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[17]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[18]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[19]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[20]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[21]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[22]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[23]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[24]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[25]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[26]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[27]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[28]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[29]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[30]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[31]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[32]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[33]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[34]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[35]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[36]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[37]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(crosslineJumpTarget_t[38]); // @[src/main/scala/nutcore/frontend/IFU.scala 334:38]
    end
    //
    if (enToggle_past) begin
      cover(r_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
  end
endmodule
module NaiveRVCAlignBuffer(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_valid, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input  [63:0] io_in_bits_instr, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input  [38:0] io_in_bits_pc, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input  [38:0] io_in_bits_pnpc, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_0, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_1, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_2, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_3, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_4, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_5, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_6, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_7, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_8, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_9, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_10, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_11, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_12, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_13, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_14, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_in_bits_exceptionVec_15, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input  [3:0]  io_in_bits_brIdx, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_out_ready, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output [63:0] io_out_bits_instr, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output [38:0] io_out_bits_pc, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output [38:0] io_out_bits_pnpc, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output        io_out_bits_exceptionVec_1, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output        io_out_bits_exceptionVec_12, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output [3:0]  io_out_bits_brIdx, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  output        io_out_bits_crossBoundaryFault, // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
  input         io_flush // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 27:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 41:22]
  wire  _instr_T = state == 2'h2; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 93:23]
  wire  _instr_T_1 = state == 2'h3; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 93:47]
  wire [79:0] instIn = {16'h0,io_in_bits_instr}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 44:19]
  reg [15:0] specialInstR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
  wire [31:0] _instr_T_4 = {instIn[15:0],specialInstR}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 93:73]
  wire  _pcOffset_T = state == 2'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 43:28]
  reg [2:0] pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 42:26]
  wire [2:0] pcOffset = state == 2'h0 ? io_in_bits_pc[2:0] : pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 43:21]
  wire  _instr_T_9 = 3'h0 == pcOffset; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _instr_T_13 = _instr_T_9 ? instIn[31:0] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _instr_T_10 = 3'h2 == pcOffset; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _instr_T_14 = _instr_T_10 ? instIn[47:16] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _instr_T_17 = _instr_T_13 | _instr_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _instr_T_11 = 3'h4 == pcOffset; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _instr_T_15 = _instr_T_11 ? instIn[63:32] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _instr_T_18 = _instr_T_17 | _instr_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _instr_T_12 = 3'h6 == pcOffset; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _instr_T_16 = _instr_T_12 ? instIn[79:48] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _instr_T_19 = _instr_T_18 | _instr_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] instr = state == 2'h2 | state == 2'h3 ? _instr_T_4 : _instr_T_19; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 93:15]
  wire  isRVC = instr[1:0] != 2'h3; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 34:27]
  wire [7:0] hasException_lo = {io_in_bits_exceptionVec_7,io_in_bits_exceptionVec_6,io_in_bits_exceptionVec_5,
    io_in_bits_exceptionVec_4,io_in_bits_exceptionVec_3,io_in_bits_exceptionVec_2,io_in_bits_exceptionVec_1,
    io_in_bits_exceptionVec_0}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 36:61]
  wire [15:0] _hasException_T = {io_in_bits_exceptionVec_15,io_in_bits_exceptionVec_14,io_in_bits_exceptionVec_13,
    io_in_bits_exceptionVec_12,io_in_bits_exceptionVec_11,io_in_bits_exceptionVec_10,io_in_bits_exceptionVec_9,
    io_in_bits_exceptionVec_8,hasException_lo}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 36:61]
  wire  hasException = io_in_valid & |_hasException_T; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 36:34]
  wire  _rvcFinish_T = pcOffset == 3'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 50:28]
  wire  _rvcFinish_T_1 = ~isRVC; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 50:40]
  wire  _rvcFinish_T_5 = pcOffset == 3'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 50:72]
  wire  _rvcFinish_T_11 = pcOffset == 3'h2; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 50:116]
  wire  _rvcFinish_T_16 = pcOffset == 3'h6; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 50:159]
  wire  rvcFinish = pcOffset == 3'h0 & (~isRVC | io_in_bits_brIdx[0]) | pcOffset == 3'h4 & (~isRVC | io_in_bits_brIdx[0]
    ) | pcOffset == 3'h2 & (isRVC | io_in_bits_brIdx[1]) | pcOffset == 3'h6 & isRVC; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 50:147]
  wire  _rvcNext_T_13 = _rvcFinish_T_11 & _rvcFinish_T_1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 53:122]
  wire  _rvcNext_T_15 = ~io_in_bits_brIdx[1]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 53:135]
  wire  rvcNext = _rvcFinish_T & (isRVC & ~io_in_bits_brIdx[0]) | _rvcFinish_T_5 & (isRVC & ~io_in_bits_brIdx[0]) |
    _rvcFinish_T_11 & _rvcFinish_T_1 & ~io_in_bits_brIdx[1]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 53:102]
  wire  _rvcSpecial_T_2 = _rvcFinish_T_16 & _rvcFinish_T_1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 54:37]
  wire  rvcSpecial = _rvcFinish_T_16 & _rvcFinish_T_1 & ~io_in_bits_brIdx[2]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 54:47]
  wire  rvcSpecialJump = _rvcSpecial_T_2 & io_in_bits_brIdx[2]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 55:51]
  wire  pnpcIsSeq = io_in_bits_brIdx[3]; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 56:24]
  wire  _flushIFU_T_2 = _pcOffset_T | state == 2'h1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 59:36]
  wire  flushIFU = (_pcOffset_T | state == 2'h1) & rvcSpecial & io_in_valid & ~pnpcIsSeq; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 59:87]
  wire  loadNextInstline = _flushIFU_T_2 & (rvcSpecial | rvcSpecialJump) & io_in_valid & pnpcIsSeq; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 62:115]
  reg [38:0] specialPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
  reg [38:0] specialNPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
  reg  specialIPFR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 69:28]
  wire  hasCrossBoundaryFault = io_in_bits_exceptionVec_1 | io_in_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 70:73]
  wire  rvcForceLoadNext = _rvcNext_T_13 & io_in_bits_pnpc[2:0] == 3'h4 & _rvcNext_T_15; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 72:86]
  wire  _canGo_T = rvcFinish | rvcNext; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 103:28]
  wire  _canIn_T = rvcFinish | rvcForceLoadNext; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 104:28]
  wire [38:0] _pnpcOut_T_1 = io_in_bits_pc + 39'h2; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 106:76]
  wire [38:0] _pnpcOut_T_3 = io_in_bits_pc + 39'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 106:95]
  wire [38:0] _pnpcOut_T_4 = isRVC ? _pnpcOut_T_1 : _pnpcOut_T_3; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 106:55]
  wire [38:0] _pnpcOut_T_5 = rvcFinish ? io_in_bits_pnpc : _pnpcOut_T_4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 106:23]
  wire  _T_6 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [1:0] _GEN_0 = _T_6 & rvcFinish ? 2'h0 : state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 107:{39,46} 41:22]
  wire [2:0] _pcOffsetR_T = isRVC ? 3'h2 : 3'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 110:38]
  wire [2:0] _pcOffsetR_T_2 = pcOffset + _pcOffsetR_T; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 110:33]
  wire [1:0] _GEN_1 = _T_6 & rvcNext ? 2'h1 : _GEN_0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 108:37 109:17]
  wire [2:0] _GEN_2 = _T_6 & rvcNext ? _pcOffsetR_T_2 : pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 108:37 110:21 42:26]
  wire [1:0] _GEN_3 = rvcSpecial & io_in_valid ? 2'h2 : _GEN_1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 112:40 113:17]
  wire [38:0] _pcOut_T_2 = {io_in_bits_pc[38:3],pcOffsetR}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 129:21]
  wire [38:0] _GEN_27 = 2'h3 == state ? specialPCR : 39'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 164:15 64:23]
  wire [38:0] _GEN_32 = 2'h2 == state ? specialPCR : _GEN_27; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 152:15]
  wire [38:0] _GEN_40 = 2'h1 == state ? _pcOut_T_2 : _GEN_32; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 129:15]
  wire [38:0] pcOut = 2'h0 == state ? io_in_bits_pc : _GEN_40; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 105:15]
  wire [38:0] _GEN_4 = rvcSpecial & io_in_valid ? pcOut : specialPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 112:40 114:22 66:23]
  wire [15:0] _GEN_5 = rvcSpecial & io_in_valid ? io_in_bits_instr[63:48] : specialInstR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 112:40 115:24 68:25]
  wire  _GEN_6 = rvcSpecial & io_in_valid ? hasCrossBoundaryFault : specialIPFR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 112:40 116:23 69:28]
  wire [1:0] _GEN_7 = rvcSpecialJump & io_in_valid ? 2'h3 : _GEN_3; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 118:44 119:17]
  wire [38:0] _GEN_8 = rvcSpecialJump & io_in_valid ? pcOut : _GEN_4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 118:44 120:22]
  wire [38:0] _GEN_9 = rvcSpecialJump & io_in_valid ? io_in_bits_pnpc : specialNPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 118:44 121:23 67:24]
  wire [15:0] _GEN_10 = rvcSpecialJump & io_in_valid ? io_in_bits_instr[63:48] : _GEN_5; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 118:44 122:24]
  wire  _GEN_11 = rvcSpecialJump & io_in_valid ? hasCrossBoundaryFault : _GEN_6; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 118:44 123:23]
  wire [38:0] _pnpcOut_T_7 = pcOut + 39'h2; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 130:68]
  wire [38:0] _pnpcOut_T_9 = pcOut + 39'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 130:79]
  wire [38:0] _pnpcOut_T_10 = isRVC ? _pnpcOut_T_7 : _pnpcOut_T_9; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 130:55]
  wire [38:0] _pnpcOut_T_11 = rvcFinish ? io_in_bits_pnpc : _pnpcOut_T_10; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 130:23]
  wire [38:0] _pnpcOut_T_13 = specialPCR + 39'h4; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 153:31]
  wire [1:0] _GEN_24 = _T_6 ? 2'h1 : state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 157:26 158:17 41:22]
  wire [2:0] _GEN_25 = _T_6 ? 3'h2 : pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 157:26 159:21 42:26]
  wire [1:0] _GEN_26 = _T_6 ? 2'h0 : state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 169:26 170:17 41:22]
  wire [38:0] _GEN_28 = 2'h3 == state ? specialNPCR : 39'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 165:17 65:25]
  wire  _GEN_29 = 2'h3 == state & io_in_valid; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 167:15 46:23]
  wire [1:0] _GEN_31 = 2'h3 == state ? _GEN_26 : state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 41:22]
  wire [38:0] _GEN_33 = 2'h2 == state ? _pnpcOut_T_13 : _GEN_28; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 153:17]
  wire  _GEN_34 = 2'h2 == state ? io_in_valid : _GEN_29; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 155:15]
  wire  _GEN_35 = 2'h2 == state ? 1'h0 : 2'h3 == state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 156:15]
  wire [1:0] _GEN_36 = 2'h2 == state ? _GEN_24 : _GEN_31; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
  wire [2:0] _GEN_37 = 2'h2 == state ? _GEN_25 : pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 42:26]
  wire  _GEN_38 = 2'h1 == state ? _canGo_T : _GEN_34; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 127:15]
  wire  _GEN_39 = 2'h1 == state ? _canIn_T : _GEN_35; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 128:15]
  wire [38:0] _GEN_41 = 2'h1 == state ? _pnpcOut_T_11 : _GEN_33; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 130:17]
  wire [1:0] _GEN_42 = 2'h1 == state ? _GEN_7 : _GEN_36; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
  wire  _GEN_48 = 2'h0 == state ? rvcFinish | rvcNext : _GEN_38; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 103:15]
  wire  canIn = 2'h0 == state ? rvcFinish | rvcForceLoadNext : _GEN_39; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 104:15]
  wire [38:0] pnpcOut = 2'h0 == state ? _pnpcOut_T_5 : _GEN_41; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 106:17]
  wire  canGo = hasException | _GEN_48; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 182:23 184:11]
  wire  _io_out_bits_brIdx_T_10 = pnpcOut == _pnpcOut_T_9 & _rvcFinish_T_1 | pnpcOut == _pnpcOut_T_7 & isRVC ? 1'h0 : 1'h1
    ; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 193:27]
  wire  _io_out_bits_exceptionVec_12_T_2 = _instr_T_1 | _instr_T; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 199:133]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [1:0] state_p; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 41:22]
  wire [1:0] state_t = state ^ state_p; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 41:22]
  wire  toggle_249_clock;
  wire  toggle_249_reset;
  wire [1:0] toggle_249_valid;
  reg [1:0] toggle_249_valid_reg;
  reg [15:0] specialInstR_p; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
  wire [15:0] specialInstR_t = specialInstR ^ specialInstR_p; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
  wire  toggle_251_clock;
  wire  toggle_251_reset;
  wire [15:0] toggle_251_valid;
  reg [15:0] toggle_251_valid_reg;
  reg [2:0] pcOffsetR_p; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 42:26]
  wire [2:0] pcOffsetR_t = pcOffsetR ^ pcOffsetR_p; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 42:26]
  wire  toggle_267_clock;
  wire  toggle_267_reset;
  wire [2:0] toggle_267_valid;
  reg [2:0] toggle_267_valid_reg;
  reg [38:0] specialPCR_p; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
  wire [38:0] specialPCR_t = specialPCR ^ specialPCR_p; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
  wire  toggle_270_clock;
  wire  toggle_270_reset;
  wire [38:0] toggle_270_valid;
  reg [38:0] toggle_270_valid_reg;
  reg [38:0] specialNPCR_p; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
  wire [38:0] specialNPCR_t = specialNPCR ^ specialNPCR_p; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
  wire  toggle_309_clock;
  wire  toggle_309_reset;
  wire [38:0] toggle_309_valid;
  reg [38:0] toggle_309_valid_reg;
  reg  specialIPFR_p; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 69:28]
  wire  specialIPFR_t = specialIPFR ^ specialIPFR_p; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 69:28]
  wire  toggle_348_clock;
  wire  toggle_348_reset;
  wire  toggle_348_valid;
  reg  toggle_348_valid_reg;
  GEN_w2_toggle #(.COVER_INDEX(249)) toggle_249 (
    .clock(toggle_249_clock),
    .reset(toggle_249_reset),
    .valid(toggle_249_valid)
  );
  GEN_w16_toggle #(.COVER_INDEX(251)) toggle_251 (
    .clock(toggle_251_clock),
    .reset(toggle_251_reset),
    .valid(toggle_251_valid)
  );
  GEN_w3_toggle #(.COVER_INDEX(267)) toggle_267 (
    .clock(toggle_267_clock),
    .reset(toggle_267_reset),
    .valid(toggle_267_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(270)) toggle_270 (
    .clock(toggle_270_clock),
    .reset(toggle_270_reset),
    .valid(toggle_270_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(309)) toggle_309 (
    .clock(toggle_309_clock),
    .reset(toggle_309_reset),
    .valid(toggle_309_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(348)) toggle_348 (
    .clock(toggle_348_clock),
    .reset(toggle_348_reset),
    .valid(toggle_348_valid)
  );
  assign io_in_ready = ~io_in_valid | _T_6 & canIn | loadNextInstline; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 196:58]
  assign io_out_valid = io_in_valid & canGo; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 195:31]
  assign io_out_bits_instr = {{32'd0}, instr}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 192:21]
  assign io_out_bits_pc = 2'h0 == state ? io_in_bits_pc : _GEN_40; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 105:15]
  assign io_out_bits_pnpc = 2'h0 == state ? _pnpcOut_T_5 : _GEN_41; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18 106:17]
  assign io_out_bits_exceptionVec_1 = io_in_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 198:28]
  assign io_out_bits_exceptionVec_12 = io_in_bits_exceptionVec_12 | specialIPFR & (_instr_T_1 | _instr_T); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 199:87]
  assign io_out_bits_brIdx = {{3'd0}, _io_out_bits_brIdx_T_10}; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 193:21]
  assign io_out_bits_crossBoundaryFault = hasCrossBoundaryFault & _io_out_bits_exceptionVec_12_T_2 & ~specialIPFR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 200:115]
  assign toggle_249_clock = clock;
  assign toggle_249_reset = reset;
  assign toggle_249_valid = state ^ toggle_249_valid_reg;
  assign toggle_251_clock = clock;
  assign toggle_251_reset = reset;
  assign toggle_251_valid = specialInstR ^ toggle_251_valid_reg;
  assign toggle_267_clock = clock;
  assign toggle_267_reset = reset;
  assign toggle_267_valid = pcOffsetR ^ toggle_267_valid_reg;
  assign toggle_270_clock = clock;
  assign toggle_270_reset = reset;
  assign toggle_270_valid = specialPCR ^ toggle_270_valid_reg;
  assign toggle_309_clock = clock;
  assign toggle_309_reset = reset;
  assign toggle_309_valid = specialNPCR ^ toggle_309_valid_reg;
  assign toggle_348_clock = clock;
  assign toggle_348_reset = reset;
  assign toggle_348_valid = specialIPFR ^ toggle_348_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 41:22]
      state <= 2'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 41:22]
    end else if (hasException) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 182:23]
      state <= 2'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 183:11]
    end else if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        state <= _GEN_7;
      end else begin
        state <= _GEN_42;
      end
    end else begin
      state <= 2'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 175:11]
    end
    if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialInstR <= _GEN_10;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialInstR <= _GEN_10;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 42:26]
      pcOffsetR <= 3'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 42:26]
    end else if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        pcOffsetR <= _GEN_2;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        pcOffsetR <= _GEN_2;
      end else begin
        pcOffsetR <= _GEN_37;
      end
    end
    if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialPCR <= _GEN_8;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialPCR <= _GEN_8;
      end
    end
    if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialNPCR <= _GEN_9;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialNPCR <= _GEN_9;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 69:28]
      specialIPFR <= 1'h0; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 69:28]
    end else if (~io_flush) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 100:18]
      if (2'h0 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialIPFR <= _GEN_11;
      end else if (2'h1 == state) begin // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 101:18]
        specialIPFR <= _GEN_11;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~flushIFU)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at NaiveIBF.scala:61 assert(!flushIFU)\n"); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 61:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    state_p <= state; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 41:22]
    toggle_249_valid_reg <= state;
    specialInstR_p <= specialInstR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
    toggle_251_valid_reg <= specialInstR;
    pcOffsetR_p <= pcOffsetR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 42:26]
    toggle_267_valid_reg <= pcOffsetR;
    specialPCR_p <= specialPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    toggle_270_valid_reg <= specialPCR;
    specialNPCR_p <= specialNPCR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    toggle_309_valid_reg <= specialNPCR;
    specialIPFR_p <= specialIPFR; // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 69:28]
    toggle_348_valid_reg <= specialIPFR;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  specialInstR = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  pcOffsetR = _RAND_2[2:0];
  _RAND_3 = {2{`RANDOM}};
  specialPCR = _RAND_3[38:0];
  _RAND_4 = {2{`RANDOM}};
  specialNPCR = _RAND_4[38:0];
  _RAND_5 = {1{`RANDOM}};
  specialIPFR = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  state_p = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  toggle_249_valid_reg = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  specialInstR_p = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  toggle_251_valid_reg = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  pcOffsetR_p = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  toggle_267_valid_reg = _RAND_11[2:0];
  _RAND_12 = {2{`RANDOM}};
  specialPCR_p = _RAND_12[38:0];
  _RAND_13 = {2{`RANDOM}};
  toggle_270_valid_reg = _RAND_13[38:0];
  _RAND_14 = {2{`RANDOM}};
  specialNPCR_p = _RAND_14[38:0];
  _RAND_15 = {2{`RANDOM}};
  toggle_309_valid_reg = _RAND_15[38:0];
  _RAND_16 = {1{`RANDOM}};
  specialIPFR_p = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  toggle_348_valid_reg = _RAND_17[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~flushIFU); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 61:9]
    end
    //
    if (enToggle_past) begin
      cover(state_t[0]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 41:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[1]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 41:22]
    end
    //
    if (enToggle_past) begin
      cover(specialInstR_t[0]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
    end
    //
    if (enToggle_past) begin
      cover(specialInstR_t[1]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
    end
    //
    if (enToggle_past) begin
      cover(specialInstR_t[2]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
    end
    //
    if (enToggle_past) begin
      cover(specialInstR_t[3]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
    end
    //
    if (enToggle_past) begin
      cover(specialInstR_t[4]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
    end
    //
    if (enToggle_past) begin
      cover(specialInstR_t[5]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
    end
    //
    if (enToggle_past) begin
      cover(specialInstR_t[6]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
    end
    //
    if (enToggle_past) begin
      cover(specialInstR_t[7]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
    end
    //
    if (enToggle_past) begin
      cover(specialInstR_t[8]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
    end
    //
    if (enToggle_past) begin
      cover(specialInstR_t[9]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
    end
    //
    if (enToggle_past) begin
      cover(specialInstR_t[10]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
    end
    //
    if (enToggle_past) begin
      cover(specialInstR_t[11]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
    end
    //
    if (enToggle_past) begin
      cover(specialInstR_t[12]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
    end
    //
    if (enToggle_past) begin
      cover(specialInstR_t[13]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
    end
    //
    if (enToggle_past) begin
      cover(specialInstR_t[14]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
    end
    //
    if (enToggle_past) begin
      cover(specialInstR_t[15]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 68:25]
    end
    //
    if (enToggle_past) begin
      cover(pcOffsetR_t[0]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 42:26]
    end
    //
    if (enToggle_past) begin
      cover(pcOffsetR_t[1]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 42:26]
    end
    //
    if (enToggle_past) begin
      cover(pcOffsetR_t[2]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 42:26]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[0]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[1]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[2]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[3]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[4]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[5]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[6]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[7]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[8]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[9]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[10]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[11]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[12]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[13]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[14]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[15]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[16]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[17]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[18]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[19]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[20]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[21]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[22]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[23]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[24]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[25]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[26]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[27]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[28]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[29]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[30]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[31]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[32]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[33]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[34]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[35]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[36]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[37]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialPCR_t[38]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 66:23]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[0]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[1]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[2]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[3]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[4]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[5]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[6]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[7]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[8]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[9]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[10]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[11]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[12]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[13]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[14]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[15]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[16]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[17]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[18]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[19]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[20]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[21]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[22]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[23]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[24]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[25]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[26]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[27]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[28]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[29]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[30]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[31]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[32]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[33]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[34]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[35]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[36]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[37]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialNPCR_t[38]); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 67:24]
    end
    //
    if (enToggle_past) begin
      cover(specialIPFR_t); // @[src/main/scala/nutcore/frontend/NaiveIBF.scala 69:28]
    end
  end
endmodule
module RVCExpander(
  input         clock,
  input         reset,
  input  [31:0] io_in, // @[src/main/scala/nutcore/frontend/RVC.scala 153:14]
  output [31:0] io_out_bits // @[src/main/scala/nutcore/frontend/RVC.scala 153:14]
);
  wire [6:0] io_out_s_opc = |io_in[12:5] ? 7'h13 : 7'h1f; // @[src/main/scala/nutcore/frontend/RVC.scala 50:20]
  wire [29:0] _io_out_s_T_7 = {io_in[10:7],io_in[12:11],io_in[5],io_in[6],2'h0,5'h2,3'h0,2'h1,io_in[4:2],io_out_s_opc}; // @[src/main/scala/nutcore/frontend/RVC.scala 51:15]
  wire [7:0] _io_out_s_T_15 = {io_in[6:5],io_in[12:10],3'h0}; // @[src/main/scala/nutcore/frontend/RVC.scala 33:18]
  wire [27:0] _io_out_s_T_20 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h7}; // @[src/main/scala/nutcore/frontend/RVC.scala 55:23]
  wire [6:0] _io_out_s_T_31 = {io_in[5],io_in[12:10],io_in[6],2'h0}; // @[src/main/scala/nutcore/frontend/RVC.scala 32:18]
  wire [26:0] _io_out_s_T_36 = {io_in[5],io_in[12:10],io_in[6],2'h0,2'h1,io_in[9:7],3'h2,2'h1,io_in[4:2],7'h3}; // @[src/main/scala/nutcore/frontend/RVC.scala 54:22]
  wire [27:0] _io_out_s_T_51 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h3}; // @[src/main/scala/nutcore/frontend/RVC.scala 53:22]
  wire [26:0] _io_out_s_T_73 = {_io_out_s_T_31[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_io_out_s_T_31[4:0],7'h3f}; // @[src/main/scala/nutcore/frontend/RVC.scala 60:25]
  wire [27:0] _io_out_s_T_93 = {_io_out_s_T_15[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_io_out_s_T_15[4:0],7'h27}; // @[src/main/scala/nutcore/frontend/RVC.scala 63:23]
  wire [26:0] _io_out_s_T_115 = {_io_out_s_T_31[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_io_out_s_T_31[4:0],7'h23}; // @[src/main/scala/nutcore/frontend/RVC.scala 62:22]
  wire [27:0] _io_out_s_T_135 = {_io_out_s_T_15[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_io_out_s_T_15[4:0],7'h23}; // @[src/main/scala/nutcore/frontend/RVC.scala 61:22]
  wire [6:0] _io_out_s_T_144 = io_in[12] ? 7'h7f : 7'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 40:25]
  wire [11:0] _io_out_s_T_146 = {_io_out_s_T_144,io_in[6:2]}; // @[src/main/scala/nutcore/frontend/RVC.scala 40:20]
  wire [31:0] io_out_s_res_8_bits = {_io_out_s_T_144,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h13}; // @[src/main/scala/nutcore/frontend/RVC.scala 72:24]
  wire  _io_out_s_opc_T_3 = |io_in[11:7]; // @[src/main/scala/nutcore/frontend/RVC.scala 74:24]
  wire [6:0] io_out_s_opc_1 = |io_in[11:7] ? 7'h1b : 7'h1f; // @[src/main/scala/nutcore/frontend/RVC.scala 74:20]
  wire [31:0] io_out_s_res_9_bits = {_io_out_s_T_144,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],io_out_s_opc_1}; // @[src/main/scala/nutcore/frontend/RVC.scala 75:15]
  wire [31:0] io_out_s_res_10_bits = {_io_out_s_T_144,io_in[6:2],5'h0,3'h0,io_in[11:7],7'h13}; // @[src/main/scala/nutcore/frontend/RVC.scala 81:22]
  wire  _io_out_s_opc_T_8 = |_io_out_s_T_146; // @[src/main/scala/nutcore/frontend/RVC.scala 87:29]
  wire [6:0] io_out_s_opc_2 = |_io_out_s_T_146 ? 7'h37 : 7'h3f; // @[src/main/scala/nutcore/frontend/RVC.scala 87:20]
  wire [14:0] _io_out_s_me_T_1 = io_in[12] ? 15'h7fff : 15'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 38:24]
  wire [31:0] _io_out_s_me_T_3 = {_io_out_s_me_T_1,io_in[6:2],12'h0}; // @[src/main/scala/nutcore/frontend/RVC.scala 38:19]
  wire [31:0] io_out_s_me_bits = {_io_out_s_me_T_3[31:12],io_in[11:7],io_out_s_opc_2}; // @[src/main/scala/nutcore/frontend/RVC.scala 88:24]
  wire [6:0] io_out_s_opc_3 = _io_out_s_opc_T_8 ? 7'h13 : 7'h1f; // @[src/main/scala/nutcore/frontend/RVC.scala 83:20]
  wire [2:0] _io_out_s_T_183 = io_in[12] ? 3'h7 : 3'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 39:29]
  wire [31:0] io_out_s_res_11_bits = {_io_out_s_T_183,io_in[4:3],io_in[5],io_in[2],io_in[6],4'h0,io_in[11:7],3'h0,io_in[
    11:7],io_out_s_opc_3}; // @[src/main/scala/nutcore/frontend/RVC.scala 84:15]
  wire [31:0] io_out_s_11_bits = io_in[11:7] == 5'h0 | io_in[11:7] == 5'h2 ? io_out_s_res_11_bits : io_out_s_me_bits; // @[src/main/scala/nutcore/frontend/RVC.scala 89:10]
  wire [25:0] _io_out_s_T_205 = {io_in[12],io_in[6:2],2'h1,io_in[9:7],3'h5,2'h1,io_in[9:7],7'h13}; // @[src/main/scala/nutcore/frontend/RVC.scala 95:21]
  wire [30:0] _GEN_0 = {{5'd0}, _io_out_s_T_205}; // @[src/main/scala/nutcore/frontend/RVC.scala 96:23]
  wire [30:0] _io_out_s_T_214 = _GEN_0 | 31'h40000000; // @[src/main/scala/nutcore/frontend/RVC.scala 96:23]
  wire [31:0] _io_out_s_T_223 = {_io_out_s_T_144,io_in[6:2],2'h1,io_in[9:7],3'h7,2'h1,io_in[9:7],7'h13}; // @[src/main/scala/nutcore/frontend/RVC.scala 97:21]
  wire [2:0] _io_out_s_funct_T_2 = {io_in[12],io_in[6:5]}; // @[src/main/scala/nutcore/frontend/RVC.scala 99:77]
  wire [30:0] io_out_s_sub = io_in[6:5] == 2'h0 ? 31'h40000000 : 31'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 100:22]
  wire [6:0] io_out_s_opc_4 = io_in[12] ? 7'h3b : 7'h33; // @[src/main/scala/nutcore/frontend/RVC.scala 101:22]
  wire [2:0] _GEN_1 = 3'h1 == _io_out_s_funct_T_2 ? 3'h4 : 3'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire [2:0] _GEN_2 = 3'h2 == _io_out_s_funct_T_2 ? 3'h6 : _GEN_1; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire [2:0] _GEN_3 = 3'h3 == _io_out_s_funct_T_2 ? 3'h7 : _GEN_2; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire [2:0] _GEN_4 = 3'h4 == _io_out_s_funct_T_2 ? 3'h0 : _GEN_3; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire [2:0] _GEN_5 = 3'h5 == _io_out_s_funct_T_2 ? 3'h0 : _GEN_4; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire [2:0] _GEN_6 = 3'h6 == _io_out_s_funct_T_2 ? 3'h2 : _GEN_5; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire [2:0] _GEN_7 = 3'h7 == _io_out_s_funct_T_2 ? 3'h3 : _GEN_6; // @[src/main/scala/nutcore/frontend/RVC.scala 102:{12,12}]
  wire [24:0] _io_out_s_T_230 = {2'h1,io_in[4:2],2'h1,io_in[9:7],_GEN_7,2'h1,io_in[9:7],io_out_s_opc_4}; // @[src/main/scala/nutcore/frontend/RVC.scala 102:12]
  wire [30:0] _GEN_8 = {{6'd0}, _io_out_s_T_230}; // @[src/main/scala/nutcore/frontend/RVC.scala 102:43]
  wire [30:0] _io_out_s_T_231 = _GEN_8 | io_out_s_sub; // @[src/main/scala/nutcore/frontend/RVC.scala 102:43]
  wire [31:0] _io_out_s_WIRE_0 = {{6'd0}, _io_out_s_T_205}; // @[src/main/scala/nutcore/frontend/RVC.scala 104:{19,19}]
  wire [31:0] _io_out_s_WIRE_1 = {{1'd0}, _io_out_s_T_214}; // @[src/main/scala/nutcore/frontend/RVC.scala 104:{19,19}]
  wire [31:0] _GEN_9 = 2'h1 == io_in[11:10] ? _io_out_s_WIRE_1 : _io_out_s_WIRE_0; // @[src/main/scala/nutcore/frontend/RVC.scala 19:{14,14}]
  wire [31:0] _GEN_10 = 2'h2 == io_in[11:10] ? _io_out_s_T_223 : _GEN_9; // @[src/main/scala/nutcore/frontend/RVC.scala 19:{14,14}]
  wire [31:0] _io_out_s_WIRE_3 = {{1'd0}, _io_out_s_T_231}; // @[src/main/scala/nutcore/frontend/RVC.scala 104:{19,19}]
  wire [31:0] io_out_s_res_12_bits = 2'h3 == io_in[11:10] ? _io_out_s_WIRE_3 : _GEN_10; // @[src/main/scala/nutcore/frontend/RVC.scala 19:{14,14}]
  wire [9:0] _io_out_s_T_241 = io_in[12] ? 10'h3ff : 10'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 41:22]
  wire [20:0] _io_out_s_T_249 = {_io_out_s_T_241,io_in[8],io_in[10:9],io_in[6],io_in[7],io_in[2],io_in[11],io_in[5:3],1'h0
    }; // @[src/main/scala/nutcore/frontend/RVC.scala 41:17]
  wire [31:0] io_out_s_res_13_bits = {_io_out_s_T_249[20],_io_out_s_T_249[10:1],_io_out_s_T_249[11],_io_out_s_T_249[19:
    12],5'h0,7'h6f}; // @[src/main/scala/nutcore/frontend/RVC.scala 91:21]
  wire [4:0] _io_out_s_T_291 = io_in[12] ? 5'h1f : 5'h0; // @[src/main/scala/nutcore/frontend/RVC.scala 42:22]
  wire [12:0] _io_out_s_T_296 = {_io_out_s_T_291,io_in[6:5],io_in[2],io_in[11:10],io_in[4:3],1'h0}; // @[src/main/scala/nutcore/frontend/RVC.scala 42:17]
  wire [31:0] io_out_s_res_14_bits = {_io_out_s_T_296[12],_io_out_s_T_296[10:5],5'h0,2'h1,io_in[9:7],3'h0,
    _io_out_s_T_296[4:1],_io_out_s_T_296[11],7'h63}; // @[src/main/scala/nutcore/frontend/RVC.scala 92:24]
  wire [31:0] io_out_s_res_15_bits = {_io_out_s_T_296[12],_io_out_s_T_296[10:5],5'h0,2'h1,io_in[9:7],3'h1,
    _io_out_s_T_296[4:1],_io_out_s_T_296[11],7'h63}; // @[src/main/scala/nutcore/frontend/RVC.scala 93:24]
  wire [6:0] io_out_s_load_opc = _io_out_s_opc_T_3 ? 7'h3 : 7'h1f; // @[src/main/scala/nutcore/frontend/RVC.scala 110:23]
  wire [25:0] _io_out_s_T_373 = {io_in[12],io_in[6:2],io_in[11:7],3'h1,io_in[11:7],7'h13}; // @[src/main/scala/nutcore/frontend/RVC.scala 111:24]
  wire [28:0] _io_out_s_T_383 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],7'h7}; // @[src/main/scala/nutcore/frontend/RVC.scala 114:25]
  wire [27:0] _io_out_s_T_392 = {io_in[3:2],io_in[12],io_in[6:4],2'h0,5'h2,3'h2,io_in[11:7],io_out_s_load_opc}; // @[src/main/scala/nutcore/frontend/RVC.scala 113:24]
  wire [28:0] _io_out_s_T_401 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],io_out_s_load_opc}; // @[src/main/scala/nutcore/frontend/RVC.scala 112:24]
  wire [19:0] _io_out_s_mv_T_2 = {io_in[6:2],3'h0,io_in[11:7],7'h13}; // @[src/main/scala/nutcore/frontend/RVC.scala 127:24]
  wire [24:0] _io_out_s_add_T_3 = {io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h33}; // @[src/main/scala/nutcore/frontend/RVC.scala 128:25]
  wire [24:0] io_out_s_jr = {io_in[6:2],io_in[11:7],3'h0,12'h67}; // @[src/main/scala/nutcore/frontend/RVC.scala 129:19]
  wire [24:0] io_out_s_reserved = {io_out_s_jr[24:7],7'h1f}; // @[src/main/scala/nutcore/frontend/RVC.scala 130:25]
  wire [24:0] _io_out_s_jr_reserved_T_2 = _io_out_s_opc_T_3 ? io_out_s_jr : io_out_s_reserved; // @[src/main/scala/nutcore/frontend/RVC.scala 131:33]
  wire  _io_out_s_jr_mv_T_1 = |io_in[6:2]; // @[src/main/scala/nutcore/frontend/RVC.scala 132:27]
  wire [31:0] io_out_s_mv_bits = {{12'd0}, _io_out_s_mv_T_2}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] io_out_s_jr_reserved_bits = {{7'd0}, _io_out_s_jr_reserved_T_2}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] io_out_s_jr_mv_bits = |io_in[6:2] ? io_out_s_mv_bits : io_out_s_jr_reserved_bits; // @[src/main/scala/nutcore/frontend/RVC.scala 132:22]
  wire [24:0] io_out_s_jalr = {io_in[6:2],io_in[11:7],3'h0,12'he7}; // @[src/main/scala/nutcore/frontend/RVC.scala 133:21]
  wire [24:0] _io_out_s_ebreak_T_1 = {io_out_s_jr[24:7],7'h73}; // @[src/main/scala/nutcore/frontend/RVC.scala 134:23]
  wire [24:0] io_out_s_ebreak = _io_out_s_ebreak_T_1 | 25'h100000; // @[src/main/scala/nutcore/frontend/RVC.scala 134:46]
  wire [24:0] _io_out_s_jalr_ebreak_T_2 = _io_out_s_opc_T_3 ? io_out_s_jalr : io_out_s_ebreak; // @[src/main/scala/nutcore/frontend/RVC.scala 135:33]
  wire [31:0] io_out_s_add_bits = {{7'd0}, _io_out_s_add_T_3}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] io_out_s_jalr_ebreak_bits = {{7'd0}, _io_out_s_jalr_ebreak_T_2}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] io_out_s_jalr_add_bits = _io_out_s_jr_mv_T_1 ? io_out_s_add_bits : io_out_s_jalr_ebreak_bits; // @[src/main/scala/nutcore/frontend/RVC.scala 136:25]
  wire [31:0] io_out_s_20_bits = io_in[12] ? io_out_s_jalr_add_bits : io_out_s_jr_mv_bits; // @[src/main/scala/nutcore/frontend/RVC.scala 137:10]
  wire [8:0] _io_out_s_T_409 = {io_in[9:7],io_in[12:10],3'h0}; // @[src/main/scala/nutcore/frontend/RVC.scala 37:20]
  wire [28:0] _io_out_s_T_416 = {_io_out_s_T_409[8:5],io_in[6:2],5'h2,3'h3,_io_out_s_T_409[4:0],7'h27}; // @[src/main/scala/nutcore/frontend/RVC.scala 121:25]
  wire [7:0] _io_out_s_T_422 = {io_in[8:7],io_in[12:9],2'h0}; // @[src/main/scala/nutcore/frontend/RVC.scala 36:20]
  wire [27:0] _io_out_s_T_429 = {_io_out_s_T_422[7:5],io_in[6:2],5'h2,3'h2,_io_out_s_T_422[4:0],7'h23}; // @[src/main/scala/nutcore/frontend/RVC.scala 120:24]
  wire [28:0] _io_out_s_T_442 = {_io_out_s_T_409[8:5],io_in[6:2],5'h2,3'h3,_io_out_s_T_409[4:0],7'h23}; // @[src/main/scala/nutcore/frontend/RVC.scala 119:24]
  wire [4:0] _io_out_T_2 = {io_in[1:0],io_in[15:13]}; // @[src/main/scala/nutcore/frontend/RVC.scala 148:10]
  wire [31:0] io_out_s_res_bits = {{2'd0}, _io_out_s_T_7}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] io_out_s_res_1_bits = {{4'd0}, _io_out_s_T_20}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_13 = 5'h1 == _io_out_T_2 ? io_out_s_res_1_bits : io_out_s_res_bits; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_2_bits = {{5'd0}, _io_out_s_T_36}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_14 = 5'h2 == _io_out_T_2 ? io_out_s_res_2_bits : _GEN_13; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_3_bits = {{4'd0}, _io_out_s_T_51}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_15 = 5'h3 == _io_out_T_2 ? io_out_s_res_3_bits : _GEN_14; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_4_bits = {{5'd0}, _io_out_s_T_73}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_16 = 5'h4 == _io_out_T_2 ? io_out_s_res_4_bits : _GEN_15; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_5_bits = {{4'd0}, _io_out_s_T_93}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_17 = 5'h5 == _io_out_T_2 ? io_out_s_res_5_bits : _GEN_16; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_6_bits = {{5'd0}, _io_out_s_T_115}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_18 = 5'h6 == _io_out_T_2 ? io_out_s_res_6_bits : _GEN_17; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_7_bits = {{4'd0}, _io_out_s_T_135}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_19 = 5'h7 == _io_out_T_2 ? io_out_s_res_7_bits : _GEN_18; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_20 = 5'h8 == _io_out_T_2 ? io_out_s_res_8_bits : _GEN_19; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_21 = 5'h9 == _io_out_T_2 ? io_out_s_res_9_bits : _GEN_20; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_22 = 5'ha == _io_out_T_2 ? io_out_s_res_10_bits : _GEN_21; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_23 = 5'hb == _io_out_T_2 ? io_out_s_11_bits : _GEN_22; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_24 = 5'hc == _io_out_T_2 ? io_out_s_res_12_bits : _GEN_23; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_25 = 5'hd == _io_out_T_2 ? io_out_s_res_13_bits : _GEN_24; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_26 = 5'he == _io_out_T_2 ? io_out_s_res_14_bits : _GEN_25; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_27 = 5'hf == _io_out_T_2 ? io_out_s_res_15_bits : _GEN_26; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_16_bits = {{6'd0}, _io_out_s_T_373}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_28 = 5'h10 == _io_out_T_2 ? io_out_s_res_16_bits : _GEN_27; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_17_bits = {{3'd0}, _io_out_s_T_383}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_29 = 5'h11 == _io_out_T_2 ? io_out_s_res_17_bits : _GEN_28; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_18_bits = {{4'd0}, _io_out_s_T_392}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_30 = 5'h12 == _io_out_T_2 ? io_out_s_res_18_bits : _GEN_29; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_19_bits = {{3'd0}, _io_out_s_T_401}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_31 = 5'h13 == _io_out_T_2 ? io_out_s_res_19_bits : _GEN_30; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_32 = 5'h14 == _io_out_T_2 ? io_out_s_20_bits : _GEN_31; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_20_bits = {{3'd0}, _io_out_s_T_416}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_33 = 5'h15 == _io_out_T_2 ? io_out_s_res_20_bits : _GEN_32; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_21_bits = {{4'd0}, _io_out_s_T_429}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_34 = 5'h16 == _io_out_T_2 ? io_out_s_res_21_bits : _GEN_33; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] io_out_s_res_22_bits = {{3'd0}, _io_out_s_T_442}; // @[src/main/scala/nutcore/frontend/RVC.scala 18:19 19:14]
  wire [31:0] _GEN_35 = 5'h17 == _io_out_T_2 ? io_out_s_res_22_bits : _GEN_34; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_36 = 5'h18 == _io_out_T_2 ? io_in : _GEN_35; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_37 = 5'h19 == _io_out_T_2 ? io_in : _GEN_36; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_38 = 5'h1a == _io_out_T_2 ? io_in : _GEN_37; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_39 = 5'h1b == _io_out_T_2 ? io_in : _GEN_38; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_40 = 5'h1c == _io_out_T_2 ? io_in : _GEN_39; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_41 = 5'h1d == _io_out_T_2 ? io_in : _GEN_40; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  wire [31:0] _GEN_42 = 5'h1e == _io_out_T_2 ? io_in : _GEN_41; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
  assign io_out_bits = 5'h1f == _io_out_T_2 ? io_in : _GEN_42; // @[src/main/scala/nutcore/frontend/RVC.scala 160:{12,12}]
endmodule
module Decoder(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_in_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [63:0] io_in_bits_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [38:0] io_in_bits_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [38:0] io_in_bits_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_in_bits_exceptionVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_in_bits_exceptionVec_12, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [3:0]  io_in_bits_brIdx, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_in_bits_crossBoundaryFault, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_out_ready, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [63:0] io_out_bits_cf_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [38:0] io_out_bits_cf_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [38:0] io_out_bits_cf_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [3:0]  io_out_bits_cf_brIdx, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_ctrl_src1Type, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_ctrl_src2Type, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [2:0]  io_out_bits_ctrl_fuType, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [6:0]  io_out_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [4:0]  io_out_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [4:0]  io_out_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_ctrl_rfWen, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [4:0]  io_out_bits_ctrl_rfDest, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_out_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output [63:0] io_out_bits_data_imm, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  output        io_isWFI, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_sfence_vma_invalid, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input         io_wfi_invalid, // @[src/main/scala/nutcore/frontend/IDU.scala 27:14]
  input  [11:0] intrVecIDU
);
  wire  expander_clock; // @[src/main/scala/nutcore/frontend/IDU.scala 35:24]
  wire  expander_reset; // @[src/main/scala/nutcore/frontend/IDU.scala 35:24]
  wire [31:0] expander_io_in; // @[src/main/scala/nutcore/frontend/IDU.scala 35:24]
  wire [31:0] expander_io_out_bits; // @[src/main/scala/nutcore/frontend/IDU.scala 35:24]
  wire [31:0] _decodeList_T = expander_io_out_bits & 32'h707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_1 = 32'h13 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_2 = expander_io_out_bits & 32'hfc00707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_3 = 32'h1013 == _decodeList_T_2; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_5 = 32'h2013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_7 = 32'h3013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_9 = 32'h4013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_11 = 32'h5013 == _decodeList_T_2; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_13 = 32'h6013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_15 = 32'h7013 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_17 = 32'h40005013 == _decodeList_T_2; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_18 = expander_io_out_bits & 32'hfe00707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_19 = 32'h33 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_21 = 32'h1033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_23 = 32'h2033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_25 = 32'h3033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_27 = 32'h4033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_29 = 32'h5033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_31 = 32'h6033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_33 = 32'h7033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_35 = 32'h40000033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_37 = 32'h40005033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_38 = expander_io_out_bits & 32'h7f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_39 = 32'h17 == _decodeList_T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_41 = 32'h37 == _decodeList_T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_43 = 32'h6f == _decodeList_T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_45 = 32'h67 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_47 = 32'h63 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_49 = 32'h1063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_51 = 32'h4063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_53 = 32'h5063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_55 = 32'h6063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_57 = 32'h7063 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_59 = 32'h3 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_61 = 32'h1003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_63 = 32'h2003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_65 = 32'h4003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_67 = 32'h5003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_69 = 32'h23 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_71 = 32'h1023 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_73 = 32'h2023 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_75 = 32'h1b == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_77 = 32'h101b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_79 = 32'h501b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_81 = 32'h4000501b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_83 = 32'h103b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_85 = 32'h503b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_87 = 32'h4000503b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_89 = 32'h3b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_91 = 32'h4000003b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_93 = 32'h6003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_95 = 32'h3003 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_97 = 32'h3023 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_99 = 32'h6b == _decodeList_T_38; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_101 = 32'h2000033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_103 = 32'h2001033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_105 = 32'h2002033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_107 = 32'h2003033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_109 = 32'h2004033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_111 = 32'h2005033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_113 = 32'h2006033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_115 = 32'h2007033 == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_117 = 32'h200003b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_119 = 32'h200403b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_121 = 32'h200503b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_123 = 32'h200603b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_125 = 32'h200703b == _decodeList_T_18; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_126 = expander_io_out_bits; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_127 = 32'h73 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_129 = 32'h100073 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_131 = 32'h30200073 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_133 = 32'hf == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_135 = 32'h10500073 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_137 = 32'h10200073 == _decodeList_T_126; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_138 = expander_io_out_bits & 32'hfe007fff; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_139 = 32'h12000073 == _decodeList_T_138; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_140 = expander_io_out_bits & 32'hf9f0707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_141 = 32'h1000302f == _decodeList_T_140; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_143 = 32'h1000202f == _decodeList_T_140; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_144 = expander_io_out_bits & 32'hf800707f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_145 = 32'h1800302f == _decodeList_T_144; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_147 = 32'h1800202f == _decodeList_T_144; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [31:0] _decodeList_T_148 = expander_io_out_bits & 32'hf800607f; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_149 = 32'h800202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_151 = 32'h202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_153 = 32'h2000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_155 = 32'h6000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_157 = 32'h4000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_159 = 32'h8000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_161 = 32'ha000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_163 = 32'hc000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_165 = 32'he000202f == _decodeList_T_148; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_167 = 32'h1073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_169 = 32'h2073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_171 = 32'h3073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_173 = 32'h5073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_175 = 32'h6073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_177 = 32'h7073 == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire  _decodeList_T_179 = 32'h100f == _decodeList_T; // @[src/main/scala/chisel3/util/Lookup.scala 31:38]
  wire [2:0] _decodeList_T_181 = _decodeList_T_177 ? 3'h4 : {{2'd0}, _decodeList_T_179}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_182 = _decodeList_T_175 ? 3'h4 : _decodeList_T_181; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_183 = _decodeList_T_173 ? 3'h4 : _decodeList_T_182; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_184 = _decodeList_T_171 ? 3'h4 : _decodeList_T_183; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_185 = _decodeList_T_169 ? 3'h4 : _decodeList_T_184; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_186 = _decodeList_T_167 ? 3'h4 : _decodeList_T_185; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_187 = _decodeList_T_165 ? 3'h5 : _decodeList_T_186; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_188 = _decodeList_T_163 ? 3'h5 : _decodeList_T_187; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_189 = _decodeList_T_161 ? 3'h5 : _decodeList_T_188; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_190 = _decodeList_T_159 ? 3'h5 : _decodeList_T_189; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_191 = _decodeList_T_157 ? 3'h5 : _decodeList_T_190; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_192 = _decodeList_T_155 ? 3'h5 : _decodeList_T_191; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_193 = _decodeList_T_153 ? 3'h5 : _decodeList_T_192; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_194 = _decodeList_T_151 ? 3'h5 : _decodeList_T_193; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_195 = _decodeList_T_149 ? 3'h5 : _decodeList_T_194; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_196 = _decodeList_T_147 ? 4'hf : {{1'd0}, _decodeList_T_195}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_197 = _decodeList_T_145 ? 4'hf : _decodeList_T_196; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_198 = _decodeList_T_143 ? 4'h5 : _decodeList_T_197; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_199 = _decodeList_T_141 ? 4'h5 : _decodeList_T_198; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_200 = _decodeList_T_139 ? 4'h5 : _decodeList_T_199; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_201 = _decodeList_T_137 ? 4'h4 : _decodeList_T_200; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_202 = _decodeList_T_135 ? 4'h4 : _decodeList_T_201; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_203 = _decodeList_T_133 ? 4'h2 : _decodeList_T_202; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_204 = _decodeList_T_131 ? 4'h4 : _decodeList_T_203; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_205 = _decodeList_T_129 ? 4'h4 : _decodeList_T_204; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_206 = _decodeList_T_127 ? 4'h4 : _decodeList_T_205; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_207 = _decodeList_T_125 ? 4'h5 : _decodeList_T_206; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_208 = _decodeList_T_123 ? 4'h5 : _decodeList_T_207; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_209 = _decodeList_T_121 ? 4'h5 : _decodeList_T_208; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_210 = _decodeList_T_119 ? 4'h5 : _decodeList_T_209; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_211 = _decodeList_T_117 ? 4'h5 : _decodeList_T_210; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_212 = _decodeList_T_115 ? 4'h5 : _decodeList_T_211; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_213 = _decodeList_T_113 ? 4'h5 : _decodeList_T_212; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_214 = _decodeList_T_111 ? 4'h5 : _decodeList_T_213; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_215 = _decodeList_T_109 ? 4'h5 : _decodeList_T_214; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_216 = _decodeList_T_107 ? 4'h5 : _decodeList_T_215; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_217 = _decodeList_T_105 ? 4'h5 : _decodeList_T_216; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_218 = _decodeList_T_103 ? 4'h5 : _decodeList_T_217; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_219 = _decodeList_T_101 ? 4'h5 : _decodeList_T_218; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_220 = _decodeList_T_99 ? 4'h4 : _decodeList_T_219; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_221 = _decodeList_T_97 ? 4'h2 : _decodeList_T_220; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_222 = _decodeList_T_95 ? 4'h4 : _decodeList_T_221; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_223 = _decodeList_T_93 ? 4'h4 : _decodeList_T_222; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_224 = _decodeList_T_91 ? 4'h5 : _decodeList_T_223; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_225 = _decodeList_T_89 ? 4'h5 : _decodeList_T_224; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_226 = _decodeList_T_87 ? 4'h5 : _decodeList_T_225; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_227 = _decodeList_T_85 ? 4'h5 : _decodeList_T_226; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_228 = _decodeList_T_83 ? 4'h5 : _decodeList_T_227; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_229 = _decodeList_T_81 ? 4'h4 : _decodeList_T_228; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_230 = _decodeList_T_79 ? 4'h4 : _decodeList_T_229; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_231 = _decodeList_T_77 ? 4'h4 : _decodeList_T_230; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_232 = _decodeList_T_75 ? 4'h4 : _decodeList_T_231; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_233 = _decodeList_T_73 ? 4'h2 : _decodeList_T_232; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_234 = _decodeList_T_71 ? 4'h2 : _decodeList_T_233; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_235 = _decodeList_T_69 ? 4'h2 : _decodeList_T_234; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_236 = _decodeList_T_67 ? 4'h4 : _decodeList_T_235; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_237 = _decodeList_T_65 ? 4'h4 : _decodeList_T_236; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_238 = _decodeList_T_63 ? 4'h4 : _decodeList_T_237; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_239 = _decodeList_T_61 ? 4'h4 : _decodeList_T_238; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_240 = _decodeList_T_59 ? 4'h4 : _decodeList_T_239; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_241 = _decodeList_T_57 ? 4'h1 : _decodeList_T_240; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_242 = _decodeList_T_55 ? 4'h1 : _decodeList_T_241; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_243 = _decodeList_T_53 ? 4'h1 : _decodeList_T_242; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_244 = _decodeList_T_51 ? 4'h1 : _decodeList_T_243; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_245 = _decodeList_T_49 ? 4'h1 : _decodeList_T_244; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_246 = _decodeList_T_47 ? 4'h1 : _decodeList_T_245; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_247 = _decodeList_T_45 ? 4'h4 : _decodeList_T_246; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_248 = _decodeList_T_43 ? 4'h7 : _decodeList_T_247; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_249 = _decodeList_T_41 ? 4'h6 : _decodeList_T_248; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_250 = _decodeList_T_39 ? 4'h6 : _decodeList_T_249; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_251 = _decodeList_T_37 ? 4'h5 : _decodeList_T_250; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_252 = _decodeList_T_35 ? 4'h5 : _decodeList_T_251; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_253 = _decodeList_T_33 ? 4'h5 : _decodeList_T_252; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_254 = _decodeList_T_31 ? 4'h5 : _decodeList_T_253; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_255 = _decodeList_T_29 ? 4'h5 : _decodeList_T_254; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_256 = _decodeList_T_27 ? 4'h5 : _decodeList_T_255; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_257 = _decodeList_T_25 ? 4'h5 : _decodeList_T_256; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_258 = _decodeList_T_23 ? 4'h5 : _decodeList_T_257; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_259 = _decodeList_T_21 ? 4'h5 : _decodeList_T_258; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_260 = _decodeList_T_19 ? 4'h5 : _decodeList_T_259; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_261 = _decodeList_T_17 ? 4'h4 : _decodeList_T_260; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_262 = _decodeList_T_15 ? 4'h4 : _decodeList_T_261; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_263 = _decodeList_T_13 ? 4'h4 : _decodeList_T_262; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_264 = _decodeList_T_11 ? 4'h4 : _decodeList_T_263; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_265 = _decodeList_T_9 ? 4'h4 : _decodeList_T_264; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_266 = _decodeList_T_7 ? 4'h4 : _decodeList_T_265; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_267 = _decodeList_T_5 ? 4'h4 : _decodeList_T_266; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] _decodeList_T_268 = _decodeList_T_3 ? 4'h4 : _decodeList_T_267; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [3:0] decodeList_0 = _decodeList_T_1 ? 4'h4 : _decodeList_T_268; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_269 = _decodeList_T_179 ? 3'h4 : 3'h3; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_270 = _decodeList_T_177 ? 3'h3 : _decodeList_T_269; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_271 = _decodeList_T_175 ? 3'h3 : _decodeList_T_270; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_272 = _decodeList_T_173 ? 3'h3 : _decodeList_T_271; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_273 = _decodeList_T_171 ? 3'h3 : _decodeList_T_272; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_274 = _decodeList_T_169 ? 3'h3 : _decodeList_T_273; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_275 = _decodeList_T_167 ? 3'h3 : _decodeList_T_274; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_276 = _decodeList_T_165 ? 3'h1 : _decodeList_T_275; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_277 = _decodeList_T_163 ? 3'h1 : _decodeList_T_276; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_278 = _decodeList_T_161 ? 3'h1 : _decodeList_T_277; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_279 = _decodeList_T_159 ? 3'h1 : _decodeList_T_278; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_280 = _decodeList_T_157 ? 3'h1 : _decodeList_T_279; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_281 = _decodeList_T_155 ? 3'h1 : _decodeList_T_280; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_282 = _decodeList_T_153 ? 3'h1 : _decodeList_T_281; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_283 = _decodeList_T_151 ? 3'h1 : _decodeList_T_282; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_284 = _decodeList_T_149 ? 3'h1 : _decodeList_T_283; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_285 = _decodeList_T_147 ? 3'h1 : _decodeList_T_284; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_286 = _decodeList_T_145 ? 3'h1 : _decodeList_T_285; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_287 = _decodeList_T_143 ? 3'h1 : _decodeList_T_286; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_288 = _decodeList_T_141 ? 3'h1 : _decodeList_T_287; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_289 = _decodeList_T_139 ? 3'h4 : _decodeList_T_288; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_290 = _decodeList_T_137 ? 3'h3 : _decodeList_T_289; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_291 = _decodeList_T_135 ? 3'h0 : _decodeList_T_290; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_292 = _decodeList_T_133 ? 3'h4 : _decodeList_T_291; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_293 = _decodeList_T_131 ? 3'h3 : _decodeList_T_292; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_294 = _decodeList_T_129 ? 3'h3 : _decodeList_T_293; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_295 = _decodeList_T_127 ? 3'h3 : _decodeList_T_294; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_296 = _decodeList_T_125 ? 3'h2 : _decodeList_T_295; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_297 = _decodeList_T_123 ? 3'h2 : _decodeList_T_296; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_298 = _decodeList_T_121 ? 3'h2 : _decodeList_T_297; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_299 = _decodeList_T_119 ? 3'h2 : _decodeList_T_298; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_300 = _decodeList_T_117 ? 3'h2 : _decodeList_T_299; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_301 = _decodeList_T_115 ? 3'h2 : _decodeList_T_300; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_302 = _decodeList_T_113 ? 3'h2 : _decodeList_T_301; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_303 = _decodeList_T_111 ? 3'h2 : _decodeList_T_302; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_304 = _decodeList_T_109 ? 3'h2 : _decodeList_T_303; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_305 = _decodeList_T_107 ? 3'h2 : _decodeList_T_304; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_306 = _decodeList_T_105 ? 3'h2 : _decodeList_T_305; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_307 = _decodeList_T_103 ? 3'h2 : _decodeList_T_306; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_308 = _decodeList_T_101 ? 3'h2 : _decodeList_T_307; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_309 = _decodeList_T_99 ? 3'h3 : _decodeList_T_308; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_310 = _decodeList_T_97 ? 3'h1 : _decodeList_T_309; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_311 = _decodeList_T_95 ? 3'h1 : _decodeList_T_310; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_312 = _decodeList_T_93 ? 3'h1 : _decodeList_T_311; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_313 = _decodeList_T_91 ? 3'h0 : _decodeList_T_312; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_314 = _decodeList_T_89 ? 3'h0 : _decodeList_T_313; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_315 = _decodeList_T_87 ? 3'h0 : _decodeList_T_314; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_316 = _decodeList_T_85 ? 3'h0 : _decodeList_T_315; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_317 = _decodeList_T_83 ? 3'h0 : _decodeList_T_316; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_318 = _decodeList_T_81 ? 3'h0 : _decodeList_T_317; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_319 = _decodeList_T_79 ? 3'h0 : _decodeList_T_318; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_320 = _decodeList_T_77 ? 3'h0 : _decodeList_T_319; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_321 = _decodeList_T_75 ? 3'h0 : _decodeList_T_320; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_322 = _decodeList_T_73 ? 3'h1 : _decodeList_T_321; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_323 = _decodeList_T_71 ? 3'h1 : _decodeList_T_322; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_324 = _decodeList_T_69 ? 3'h1 : _decodeList_T_323; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_325 = _decodeList_T_67 ? 3'h1 : _decodeList_T_324; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_326 = _decodeList_T_65 ? 3'h1 : _decodeList_T_325; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_327 = _decodeList_T_63 ? 3'h1 : _decodeList_T_326; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_328 = _decodeList_T_61 ? 3'h1 : _decodeList_T_327; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_329 = _decodeList_T_59 ? 3'h1 : _decodeList_T_328; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_330 = _decodeList_T_57 ? 3'h0 : _decodeList_T_329; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_331 = _decodeList_T_55 ? 3'h0 : _decodeList_T_330; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_332 = _decodeList_T_53 ? 3'h0 : _decodeList_T_331; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_333 = _decodeList_T_51 ? 3'h0 : _decodeList_T_332; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_334 = _decodeList_T_49 ? 3'h0 : _decodeList_T_333; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_335 = _decodeList_T_47 ? 3'h0 : _decodeList_T_334; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_336 = _decodeList_T_45 ? 3'h0 : _decodeList_T_335; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_337 = _decodeList_T_43 ? 3'h0 : _decodeList_T_336; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_338 = _decodeList_T_41 ? 3'h0 : _decodeList_T_337; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_339 = _decodeList_T_39 ? 3'h0 : _decodeList_T_338; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_340 = _decodeList_T_37 ? 3'h0 : _decodeList_T_339; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_341 = _decodeList_T_35 ? 3'h0 : _decodeList_T_340; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_342 = _decodeList_T_33 ? 3'h0 : _decodeList_T_341; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_343 = _decodeList_T_31 ? 3'h0 : _decodeList_T_342; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_344 = _decodeList_T_29 ? 3'h0 : _decodeList_T_343; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_345 = _decodeList_T_27 ? 3'h0 : _decodeList_T_344; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_346 = _decodeList_T_25 ? 3'h0 : _decodeList_T_345; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_347 = _decodeList_T_23 ? 3'h0 : _decodeList_T_346; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_348 = _decodeList_T_21 ? 3'h0 : _decodeList_T_347; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_349 = _decodeList_T_19 ? 3'h0 : _decodeList_T_348; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_350 = _decodeList_T_17 ? 3'h0 : _decodeList_T_349; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_351 = _decodeList_T_15 ? 3'h0 : _decodeList_T_350; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_352 = _decodeList_T_13 ? 3'h0 : _decodeList_T_351; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_353 = _decodeList_T_11 ? 3'h0 : _decodeList_T_352; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_354 = _decodeList_T_9 ? 3'h0 : _decodeList_T_353; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_355 = _decodeList_T_7 ? 3'h0 : _decodeList_T_354; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_356 = _decodeList_T_5 ? 3'h0 : _decodeList_T_355; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_357 = _decodeList_T_3 ? 3'h0 : _decodeList_T_356; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] decodeList_1 = _decodeList_T_1 ? 3'h0 : _decodeList_T_357; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_359 = _decodeList_T_177 ? 3'h7 : {{2'd0}, _decodeList_T_179}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_360 = _decodeList_T_175 ? 3'h6 : _decodeList_T_359; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_361 = _decodeList_T_173 ? 3'h5 : _decodeList_T_360; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_362 = _decodeList_T_171 ? 3'h3 : _decodeList_T_361; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_363 = _decodeList_T_169 ? 3'h2 : _decodeList_T_362; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [2:0] _decodeList_T_364 = _decodeList_T_167 ? 3'h1 : _decodeList_T_363; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_365 = _decodeList_T_165 ? 6'h32 : {{3'd0}, _decodeList_T_364}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_366 = _decodeList_T_163 ? 6'h31 : _decodeList_T_365; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_367 = _decodeList_T_161 ? 6'h30 : _decodeList_T_366; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_368 = _decodeList_T_159 ? 6'h37 : _decodeList_T_367; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_369 = _decodeList_T_157 ? 6'h26 : _decodeList_T_368; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_370 = _decodeList_T_155 ? 6'h25 : _decodeList_T_369; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [5:0] _decodeList_T_371 = _decodeList_T_153 ? 6'h24 : _decodeList_T_370; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_372 = _decodeList_T_151 ? 7'h63 : {{1'd0}, _decodeList_T_371}; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_373 = _decodeList_T_149 ? 7'h22 : _decodeList_T_372; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_374 = _decodeList_T_147 ? 7'h21 : _decodeList_T_373; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_375 = _decodeList_T_145 ? 7'h21 : _decodeList_T_374; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_376 = _decodeList_T_143 ? 7'h20 : _decodeList_T_375; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_377 = _decodeList_T_141 ? 7'h20 : _decodeList_T_376; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_378 = _decodeList_T_139 ? 7'h2 : _decodeList_T_377; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_379 = _decodeList_T_137 ? 7'h0 : _decodeList_T_378; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_380 = _decodeList_T_135 ? 7'h40 : _decodeList_T_379; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_381 = _decodeList_T_133 ? 7'h0 : _decodeList_T_380; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_382 = _decodeList_T_131 ? 7'h0 : _decodeList_T_381; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_383 = _decodeList_T_129 ? 7'h0 : _decodeList_T_382; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_384 = _decodeList_T_127 ? 7'h0 : _decodeList_T_383; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_385 = _decodeList_T_125 ? 7'hf : _decodeList_T_384; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_386 = _decodeList_T_123 ? 7'he : _decodeList_T_385; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_387 = _decodeList_T_121 ? 7'hd : _decodeList_T_386; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_388 = _decodeList_T_119 ? 7'hc : _decodeList_T_387; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_389 = _decodeList_T_117 ? 7'h8 : _decodeList_T_388; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_390 = _decodeList_T_115 ? 7'h7 : _decodeList_T_389; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_391 = _decodeList_T_113 ? 7'h6 : _decodeList_T_390; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_392 = _decodeList_T_111 ? 7'h5 : _decodeList_T_391; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_393 = _decodeList_T_109 ? 7'h4 : _decodeList_T_392; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_394 = _decodeList_T_107 ? 7'h3 : _decodeList_T_393; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_395 = _decodeList_T_105 ? 7'h2 : _decodeList_T_394; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_396 = _decodeList_T_103 ? 7'h1 : _decodeList_T_395; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_397 = _decodeList_T_101 ? 7'h0 : _decodeList_T_396; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_398 = _decodeList_T_99 ? 7'h2 : _decodeList_T_397; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_399 = _decodeList_T_97 ? 7'hb : _decodeList_T_398; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_400 = _decodeList_T_95 ? 7'h3 : _decodeList_T_399; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_401 = _decodeList_T_93 ? 7'h6 : _decodeList_T_400; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_402 = _decodeList_T_91 ? 7'h28 : _decodeList_T_401; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_403 = _decodeList_T_89 ? 7'h60 : _decodeList_T_402; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_404 = _decodeList_T_87 ? 7'h2d : _decodeList_T_403; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_405 = _decodeList_T_85 ? 7'h25 : _decodeList_T_404; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_406 = _decodeList_T_83 ? 7'h21 : _decodeList_T_405; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_407 = _decodeList_T_81 ? 7'h2d : _decodeList_T_406; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_408 = _decodeList_T_79 ? 7'h25 : _decodeList_T_407; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_409 = _decodeList_T_77 ? 7'h21 : _decodeList_T_408; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_410 = _decodeList_T_75 ? 7'h60 : _decodeList_T_409; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_411 = _decodeList_T_73 ? 7'ha : _decodeList_T_410; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_412 = _decodeList_T_71 ? 7'h9 : _decodeList_T_411; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_413 = _decodeList_T_69 ? 7'h8 : _decodeList_T_412; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_414 = _decodeList_T_67 ? 7'h5 : _decodeList_T_413; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_415 = _decodeList_T_65 ? 7'h4 : _decodeList_T_414; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_416 = _decodeList_T_63 ? 7'h2 : _decodeList_T_415; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_417 = _decodeList_T_61 ? 7'h1 : _decodeList_T_416; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_418 = _decodeList_T_59 ? 7'h0 : _decodeList_T_417; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_419 = _decodeList_T_57 ? 7'h17 : _decodeList_T_418; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_420 = _decodeList_T_55 ? 7'h16 : _decodeList_T_419; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_421 = _decodeList_T_53 ? 7'h15 : _decodeList_T_420; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_422 = _decodeList_T_51 ? 7'h14 : _decodeList_T_421; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_423 = _decodeList_T_49 ? 7'h11 : _decodeList_T_422; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_424 = _decodeList_T_47 ? 7'h10 : _decodeList_T_423; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_425 = _decodeList_T_45 ? 7'h5a : _decodeList_T_424; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_426 = _decodeList_T_43 ? 7'h58 : _decodeList_T_425; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_427 = _decodeList_T_41 ? 7'h40 : _decodeList_T_426; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_428 = _decodeList_T_39 ? 7'h40 : _decodeList_T_427; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_429 = _decodeList_T_37 ? 7'hd : _decodeList_T_428; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_430 = _decodeList_T_35 ? 7'h8 : _decodeList_T_429; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_431 = _decodeList_T_33 ? 7'h7 : _decodeList_T_430; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_432 = _decodeList_T_31 ? 7'h6 : _decodeList_T_431; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_433 = _decodeList_T_29 ? 7'h5 : _decodeList_T_432; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_434 = _decodeList_T_27 ? 7'h4 : _decodeList_T_433; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_435 = _decodeList_T_25 ? 7'h3 : _decodeList_T_434; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_436 = _decodeList_T_23 ? 7'h2 : _decodeList_T_435; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_437 = _decodeList_T_21 ? 7'h1 : _decodeList_T_436; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_438 = _decodeList_T_19 ? 7'h40 : _decodeList_T_437; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_439 = _decodeList_T_17 ? 7'hd : _decodeList_T_438; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_440 = _decodeList_T_15 ? 7'h7 : _decodeList_T_439; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_441 = _decodeList_T_13 ? 7'h6 : _decodeList_T_440; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_442 = _decodeList_T_11 ? 7'h5 : _decodeList_T_441; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_443 = _decodeList_T_9 ? 7'h4 : _decodeList_T_442; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_444 = _decodeList_T_7 ? 7'h3 : _decodeList_T_443; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_445 = _decodeList_T_5 ? 7'h2 : _decodeList_T_444; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] _decodeList_T_446 = _decodeList_T_3 ? 7'h1 : _decodeList_T_445; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire [6:0] decodeList_2 = _decodeList_T_1 ? 7'h40 : _decodeList_T_446; // @[src/main/scala/chisel3/util/Lookup.scala 34:39]
  wire  hasIntr = |intrVecIDU; // @[src/main/scala/nutcore/frontend/IDU.scala 130:22]
  wire [3:0] instrType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 4'h0 : decodeList_0; // @[src/main/scala/nutcore/frontend/IDU.scala 45:75]
  wire [2:0] fuType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 3'h3 : decodeList_1; // @[src/main/scala/nutcore/frontend/IDU.scala 45:75]
  wire [6:0] fuOpType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 7'h0 : decodeList_2; // @[src/main/scala/nutcore/frontend/IDU.scala 45:75]
  wire  _src1Type_T = 4'h4 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_2 = 4'h2 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_3 = 4'hf == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_4 = 4'h1 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_5 = 4'h6 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_6 = 4'h7 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _src1Type_T_7 = 4'h0 == instrType; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  src1Type = _src1Type_T_5 | _src1Type_T_6 | _src1Type_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  src2Type = _src1Type_T | _src1Type_T_5 | _src1Type_T_6 | _src1Type_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [4:0] rs = expander_io_out_bits[19:15]; // @[src/main/scala/nutcore/frontend/IDU.scala 65:28]
  wire [4:0] rt = expander_io_out_bits[24:20]; // @[src/main/scala/nutcore/frontend/IDU.scala 65:43]
  wire [4:0] rd = expander_io_out_bits[11:7]; // @[src/main/scala/nutcore/frontend/IDU.scala 65:58]
  wire  imm_signBit = expander_io_out_bits[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [51:0] _imm_T_1 = imm_signBit ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imm_T_2 = {_imm_T_1,expander_io_out_bits[31:20]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [11:0] _imm_T_5 = {expander_io_out_bits[31:25],rd}; // @[src/main/scala/nutcore/frontend/IDU.scala 82:27]
  wire  imm_signBit_1 = _imm_T_5[11]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [51:0] _imm_T_6 = imm_signBit_1 ? 52'hfffffffffffff : 52'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imm_T_7 = {_imm_T_6,expander_io_out_bits[31:25],rd}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [12:0] _imm_T_17 = {expander_io_out_bits[31],expander_io_out_bits[7],expander_io_out_bits[30:25],
    expander_io_out_bits[11:8],1'h0}; // @[src/main/scala/nutcore/frontend/IDU.scala 84:27]
  wire  imm_signBit_3 = _imm_T_17[12]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [50:0] _imm_T_18 = imm_signBit_3 ? 51'h7ffffffffffff : 51'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imm_T_19 = {_imm_T_18,expander_io_out_bits[31],expander_io_out_bits[7],expander_io_out_bits[30:25],
    expander_io_out_bits[11:8],1'h0}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [31:0] _imm_T_21 = {expander_io_out_bits[31:12],12'h0}; // @[src/main/scala/nutcore/frontend/IDU.scala 85:27]
  wire  imm_signBit_4 = _imm_T_21[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _imm_T_22 = imm_signBit_4 ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imm_T_23 = {_imm_T_22,expander_io_out_bits[31:12],12'h0}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [20:0] _imm_T_28 = {expander_io_out_bits[31],expander_io_out_bits[19:12],expander_io_out_bits[20],
    expander_io_out_bits[30:21],1'h0}; // @[src/main/scala/nutcore/frontend/IDU.scala 86:27]
  wire  imm_signBit_5 = _imm_T_28[20]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [42:0] _imm_T_29 = imm_signBit_5 ? 43'h7ffffffffff : 43'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imm_T_30 = {_imm_T_29,expander_io_out_bits[31],expander_io_out_bits[19:12],expander_io_out_bits[20],
    expander_io_out_bits[30:21],1'h0}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _imm_T_37 = _src1Type_T ? _imm_T_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_38 = _src1Type_T_2 ? _imm_T_7 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_39 = _src1Type_T_3 ? _imm_T_7 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_40 = _src1Type_T_4 ? _imm_T_19 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_41 = _src1Type_T_5 ? _imm_T_23 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_42 = _src1Type_T_6 ? _imm_T_30 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_43 = _imm_T_37 | _imm_T_38; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_44 = _imm_T_43 | _imm_T_39; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_45 = _imm_T_44 | _imm_T_40; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _imm_T_46 = _imm_T_45 | _imm_T_41; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _T_9 = rd == 5'h1 | rd == 5'h5; // @[src/main/scala/nutcore/frontend/IDU.scala 91:42]
  wire [6:0] _GEN_0 = _T_9 & fuOpType == 7'h58 ? 7'h5c : fuOpType; // @[src/main/scala/nutcore/frontend/IDU.scala 50:29 92:{57,85}]
  wire  _T_15 = rs == 5'h1 | rs == 5'h5; // @[src/main/scala/nutcore/frontend/IDU.scala 91:42]
  wire [6:0] _GEN_1 = _T_15 ? 7'h5e : _GEN_0; // @[src/main/scala/nutcore/frontend/IDU.scala 94:{29,57}]
  wire [6:0] _GEN_2 = _T_9 ? 7'h5c : _GEN_1; // @[src/main/scala/nutcore/frontend/IDU.scala 95:{29,57}]
  wire [6:0] _GEN_3 = fuOpType == 7'h5a ? _GEN_2 : _GEN_0; // @[src/main/scala/nutcore/frontend/IDU.scala 93:40]
  wire  _io_in_ready_T_1 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  is_sfence_vma = fuType == 3'h4 & fuOpType == 7'h2; // @[src/main/scala/nutcore/frontend/IDU.scala 136:45]
  wire  sfence_vma_illegal = is_sfence_vma & io_sfence_vma_invalid; // @[src/main/scala/nutcore/frontend/IDU.scala 137:42]
  wire  wfi_illegal = io_isWFI & io_wfi_invalid; // @[src/main/scala/nutcore/frontend/IDU.scala 138:30]
  wire  illegal_instr = instrType == 4'h0 | sfence_vma_illegal | wfi_illegal; // @[src/main/scala/nutcore/frontend/IDU.scala 139:82]
  RVCExpander expander ( // @[src/main/scala/nutcore/frontend/IDU.scala 35:24]
    .clock(expander_clock),
    .reset(expander_reset),
    .io_in(expander_io_in),
    .io_out_bits(expander_io_out_bits)
  );
  assign io_in_ready = ~io_in_valid | _io_in_ready_T_1; // @[src/main/scala/nutcore/frontend/IDU.scala 120:31]
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 119:16]
  assign io_out_bits_cf_instr = io_in_bits_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 121:18]
  assign io_out_bits_cf_pc = io_in_bits_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 121:18]
  assign io_out_bits_cf_pnpc = io_in_bits_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 121:18]
  assign io_out_bits_cf_exceptionVec_1 = io_in_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 142:49]
  assign io_out_bits_cf_exceptionVec_2 = illegal_instr & ~hasIntr & io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 140:74]
  assign io_out_bits_cf_exceptionVec_12 = io_in_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/IDU.scala 141:47]
  assign io_out_bits_cf_intrVec_1 = intrVecIDU[1]; // @[src/main/scala/nutcore/frontend/IDU.scala 129:38]
  assign io_out_bits_cf_intrVec_3 = intrVecIDU[3]; // @[src/main/scala/nutcore/frontend/IDU.scala 129:38]
  assign io_out_bits_cf_intrVec_5 = intrVecIDU[5]; // @[src/main/scala/nutcore/frontend/IDU.scala 129:38]
  assign io_out_bits_cf_intrVec_7 = intrVecIDU[7]; // @[src/main/scala/nutcore/frontend/IDU.scala 129:38]
  assign io_out_bits_cf_intrVec_9 = intrVecIDU[9]; // @[src/main/scala/nutcore/frontend/IDU.scala 129:38]
  assign io_out_bits_cf_intrVec_11 = intrVecIDU[11]; // @[src/main/scala/nutcore/frontend/IDU.scala 129:38]
  assign io_out_bits_cf_brIdx = io_in_bits_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 121:18]
  assign io_out_bits_cf_crossBoundaryFault = io_in_bits_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/IDU.scala 121:18]
  assign io_out_bits_ctrl_src1Type = expander_io_out_bits[6:0] == 7'h37 ? 1'h0 : src1Type; // @[src/main/scala/nutcore/frontend/IDU.scala 99:35]
  assign io_out_bits_ctrl_src2Type = _src1Type_T | _src1Type_T_5 | _src1Type_T_6 | _src1Type_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_bits_ctrl_fuType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 3'h3 :
    decodeList_1; // @[src/main/scala/nutcore/frontend/IDU.scala 45:75]
  assign io_out_bits_ctrl_fuOpType = fuType == 3'h0 ? _GEN_3 : fuOpType; // @[src/main/scala/nutcore/frontend/IDU.scala 50:29 90:32]
  assign io_out_bits_ctrl_rfSrc1 = src1Type ? 5'h0 : rs; // @[src/main/scala/nutcore/frontend/IDU.scala 74:33]
  assign io_out_bits_ctrl_rfSrc2 = ~src2Type ? rt : 5'h0; // @[src/main/scala/nutcore/frontend/IDU.scala 75:33]
  assign io_out_bits_ctrl_rfWen = instrType[2]; // @[src/main/scala/nutcore/Decode.scala 33:50]
  assign io_out_bits_ctrl_rfDest = instrType[2] ? rd : 5'h0; // @[src/main/scala/nutcore/frontend/IDU.scala 77:33]
  assign io_out_bits_ctrl_isNutCoreTrap = _decodeList_T_99 & io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 144:66]
  assign io_out_bits_data_imm = _imm_T_46 | _imm_T_42; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_isWFI = _decodeList_T_135 & io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 145:43]
  assign expander_clock = clock;
  assign expander_reset = reset;
  assign expander_io_in = io_in_bits_instr[31:0]; // @[src/main/scala/nutcore/frontend/IDU.scala 36:18]
endmodule
module IDU(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_in_0_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input  [63:0] io_in_0_bits_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input  [38:0] io_in_0_bits_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input  [38:0] io_in_0_bits_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_in_0_bits_exceptionVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_in_0_bits_exceptionVec_12, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input  [3:0]  io_in_0_bits_brIdx, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_in_0_bits_crossBoundaryFault, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_out_0_ready, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_valid, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [63:0] io_out_0_bits_cf_instr, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [38:0] io_out_0_bits_cf_pc, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [38:0] io_out_0_bits_cf_pnpc, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [3:0]  io_out_0_bits_cf_brIdx, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_ctrl_src1Type, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_ctrl_src2Type, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [2:0]  io_out_0_bits_ctrl_fuType, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [6:0]  io_out_0_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [4:0]  io_out_0_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [4:0]  io_out_0_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_ctrl_rfWen, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [4:0]  io_out_0_bits_ctrl_rfDest, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        io_out_0_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output [63:0] io_out_0_bits_data_imm, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_sfence_vma_invalid, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  input         io_wfi_invalid, // @[src/main/scala/nutcore/frontend/IDU.scala 164:14]
  output        isWFI_0,
  input  [11:0] intrVecIDU
);
  wire  decoder_clock; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_reset; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_in_ready; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_in_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [63:0] decoder_io_in_bits_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [38:0] decoder_io_in_bits_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [38:0] decoder_io_in_bits_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_in_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_in_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [3:0] decoder_io_in_bits_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_in_bits_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_ready; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [63:0] decoder_io_out_bits_cf_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [38:0] decoder_io_out_bits_cf_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [38:0] decoder_io_out_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [3:0] decoder_io_out_bits_cf_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_ctrl_src1Type; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_ctrl_src2Type; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [2:0] decoder_io_out_bits_ctrl_fuType; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [6:0] decoder_io_out_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [4:0] decoder_io_out_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [4:0] decoder_io_out_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_ctrl_rfWen; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [4:0] decoder_io_out_bits_ctrl_rfDest; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_out_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [63:0] decoder_io_out_bits_data_imm; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_isWFI; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_sfence_vma_invalid; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  decoder_io_wfi_invalid; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire [11:0] decoder_intrVecIDU; // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
  wire  isWFI = decoder_io_isWFI; // @[src/main/scala/nutcore/frontend/IDU.scala 175:{23,23}]
  Decoder decoder ( // @[src/main/scala/nutcore/frontend/IDU.scala 170:23]
    .clock(decoder_clock),
    .reset(decoder_reset),
    .io_in_ready(decoder_io_in_ready),
    .io_in_valid(decoder_io_in_valid),
    .io_in_bits_instr(decoder_io_in_bits_instr),
    .io_in_bits_pc(decoder_io_in_bits_pc),
    .io_in_bits_pnpc(decoder_io_in_bits_pnpc),
    .io_in_bits_exceptionVec_1(decoder_io_in_bits_exceptionVec_1),
    .io_in_bits_exceptionVec_12(decoder_io_in_bits_exceptionVec_12),
    .io_in_bits_brIdx(decoder_io_in_bits_brIdx),
    .io_in_bits_crossBoundaryFault(decoder_io_in_bits_crossBoundaryFault),
    .io_out_ready(decoder_io_out_ready),
    .io_out_valid(decoder_io_out_valid),
    .io_out_bits_cf_instr(decoder_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(decoder_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(decoder_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(decoder_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(decoder_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_exceptionVec_12(decoder_io_out_bits_cf_exceptionVec_12),
    .io_out_bits_cf_intrVec_1(decoder_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_3(decoder_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_5(decoder_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_7(decoder_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_9(decoder_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_11(decoder_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(decoder_io_out_bits_cf_brIdx),
    .io_out_bits_cf_crossBoundaryFault(decoder_io_out_bits_cf_crossBoundaryFault),
    .io_out_bits_ctrl_src1Type(decoder_io_out_bits_ctrl_src1Type),
    .io_out_bits_ctrl_src2Type(decoder_io_out_bits_ctrl_src2Type),
    .io_out_bits_ctrl_fuType(decoder_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(decoder_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_rfSrc1(decoder_io_out_bits_ctrl_rfSrc1),
    .io_out_bits_ctrl_rfSrc2(decoder_io_out_bits_ctrl_rfSrc2),
    .io_out_bits_ctrl_rfWen(decoder_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(decoder_io_out_bits_ctrl_rfDest),
    .io_out_bits_ctrl_isNutCoreTrap(decoder_io_out_bits_ctrl_isNutCoreTrap),
    .io_out_bits_data_imm(decoder_io_out_bits_data_imm),
    .io_isWFI(decoder_io_isWFI),
    .io_sfence_vma_invalid(decoder_io_sfence_vma_invalid),
    .io_wfi_invalid(decoder_io_wfi_invalid),
    .intrVecIDU(decoder_intrVecIDU)
  );
  assign io_in_0_ready = decoder_io_in_ready; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign io_out_0_valid = decoder_io_out_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_instr = decoder_io_out_bits_cf_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_pc = decoder_io_out_bits_cf_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_pnpc = decoder_io_out_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_exceptionVec_1 = decoder_io_out_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_exceptionVec_2 = decoder_io_out_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_exceptionVec_12 = decoder_io_out_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_intrVec_1 = decoder_io_out_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_intrVec_3 = decoder_io_out_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_intrVec_5 = decoder_io_out_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_intrVec_7 = decoder_io_out_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_intrVec_9 = decoder_io_out_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_intrVec_11 = decoder_io_out_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_brIdx = decoder_io_out_bits_cf_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_cf_crossBoundaryFault = decoder_io_out_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_src1Type = decoder_io_out_bits_ctrl_src1Type; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_src2Type = decoder_io_out_bits_ctrl_src2Type; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_fuType = decoder_io_out_bits_ctrl_fuType; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_fuOpType = decoder_io_out_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_rfSrc1 = decoder_io_out_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_rfSrc2 = decoder_io_out_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_rfWen = decoder_io_out_bits_ctrl_rfWen; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_rfDest = decoder_io_out_bits_ctrl_rfDest; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_ctrl_isNutCoreTrap = decoder_io_out_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign io_out_0_bits_data_imm = decoder_io_out_bits_data_imm; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign isWFI_0 = isWFI;
  assign decoder_clock = clock;
  assign decoder_reset = reset;
  assign decoder_io_in_valid = io_in_0_valid; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_instr = io_in_0_bits_instr; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_pc = io_in_0_bits_pc; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_pnpc = io_in_0_bits_pnpc; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_exceptionVec_1 = io_in_0_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_exceptionVec_12 = io_in_0_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_brIdx = io_in_0_bits_brIdx; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_in_bits_crossBoundaryFault = io_in_0_bits_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/IDU.scala 173:12]
  assign decoder_io_out_ready = io_out_0_ready; // @[src/main/scala/nutcore/frontend/IDU.scala 174:13]
  assign decoder_io_sfence_vma_invalid = io_sfence_vma_invalid; // @[src/main/scala/nutcore/frontend/IDU.scala 171:33]
  assign decoder_io_wfi_invalid = io_wfi_invalid; // @[src/main/scala/nutcore/frontend/IDU.scala 172:26]
  assign decoder_intrVecIDU = intrVecIDU;
endmodule
module FlushableQueue(
  input         clock,
  input         reset,
  output        io_enq_ready, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input         io_enq_valid, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input  [63:0] io_enq_bits_instr, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input  [38:0] io_enq_bits_pc, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input  [38:0] io_enq_bits_pnpc, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input         io_enq_bits_exceptionVec_1, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input  [3:0]  io_enq_bits_brIdx, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input         io_deq_ready, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_valid, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output [63:0] io_deq_bits_instr, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output [38:0] io_deq_bits_pc, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output [38:0] io_deq_bits_pnpc, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_0, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_1, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_2, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_3, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_4, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_5, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_6, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_7, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_8, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_9, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_10, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_11, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_12, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_13, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_14, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output        io_deq_bits_exceptionVec_15, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  output [3:0]  io_deq_bits_brIdx, // @[src/main/scala/utils/FlushableQueue.scala 21:14]
  input         io_flush // @[src/main/scala/utils/FlushableQueue.scala 21:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_instr [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_instr_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_instr_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [63:0] ram_instr_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [63:0] ram_instr_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_instr_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_instr_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_instr_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg [38:0] ram_pc [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pc_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_pc_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [38:0] ram_pc_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [38:0] ram_pc_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_pc_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pc_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pc_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg [38:0] ram_pnpc [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pnpc_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_pnpc_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [38:0] ram_pnpc_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [38:0] ram_pnpc_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_pnpc_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pnpc_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_pnpc_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_0 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_0_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_0_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_0_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_0_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_0_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_0_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_0_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_1 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_1_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_1_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_1_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_1_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_1_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_1_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_1_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_2 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_2_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_2_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_2_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_2_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_2_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_2_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_2_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_3 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_3_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_3_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_3_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_3_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_3_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_3_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_3_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_4 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_4_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_4_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_4_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_4_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_4_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_4_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_4_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_5 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_5_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_5_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_5_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_5_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_5_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_5_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_5_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_6 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_6_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_6_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_6_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_6_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_6_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_6_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_6_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_7 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_7_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_7_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_7_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_7_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_7_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_7_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_7_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_8 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_8_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_8_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_8_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_8_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_8_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_8_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_8_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_9 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_9_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_9_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_9_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_9_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_9_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_9_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_9_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_10 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_10_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_10_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_10_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_10_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_10_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_10_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_10_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_11 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_11_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_11_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_11_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_11_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_11_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_11_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_11_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_12 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_12_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_12_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_12_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_12_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_12_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_12_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_12_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_13 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_13_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_13_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_13_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_13_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_13_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_13_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_13_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_14 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_14_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_14_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_14_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_14_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_14_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_14_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_14_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg  ram_exceptionVec_15 [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_15_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_15_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_15_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_15_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_exceptionVec_15_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_15_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_exceptionVec_15_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg [3:0] ram_brIdx [0:3]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_brIdx_io_deq_bits_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_brIdx_io_deq_bits_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [3:0] ram_brIdx_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [3:0] ram_brIdx_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire [1:0] ram_brIdx_MPORT_addr; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_brIdx_MPORT_mask; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  wire  ram_brIdx_MPORT_en; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  reg [1:0] enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  maybe_full; // @[src/main/scala/utils/FlushableQueue.scala 26:35]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[src/main/scala/utils/FlushableQueue.scala 28:41]
  wire  empty = ptr_match & ~maybe_full; // @[src/main/scala/utils/FlushableQueue.scala 29:33]
  wire  full = ptr_match & maybe_full; // @[src/main/scala/utils/FlushableQueue.scala 30:32]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [1:0] enq_ptr_value_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [1:0] enq_ptr_value_t = enq_ptr_value ^ enq_ptr_value_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  toggle_349_clock;
  wire  toggle_349_reset;
  wire [1:0] toggle_349_valid;
  reg [1:0] toggle_349_valid_reg;
  reg [1:0] deq_ptr_value_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [1:0] deq_ptr_value_t = deq_ptr_value ^ deq_ptr_value_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  toggle_351_clock;
  wire  toggle_351_reset;
  wire [1:0] toggle_351_valid;
  reg [1:0] toggle_351_valid_reg;
  reg  maybe_full_p; // @[src/main/scala/utils/FlushableQueue.scala 26:35]
  wire  maybe_full_t = maybe_full ^ maybe_full_p; // @[src/main/scala/utils/FlushableQueue.scala 26:35]
  wire  toggle_353_clock;
  wire  toggle_353_reset;
  wire  toggle_353_valid;
  reg  toggle_353_valid_reg;
  GEN_w2_toggle #(.COVER_INDEX(349)) toggle_349 (
    .clock(toggle_349_clock),
    .reset(toggle_349_reset),
    .valid(toggle_349_valid)
  );
  GEN_w2_toggle #(.COVER_INDEX(351)) toggle_351 (
    .clock(toggle_351_clock),
    .reset(toggle_351_reset),
    .valid(toggle_351_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(353)) toggle_353 (
    .clock(toggle_353_clock),
    .reset(toggle_353_reset),
    .valid(toggle_353_valid)
  );
  assign ram_instr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_instr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_instr_io_deq_bits_MPORT_data = ram_instr[ram_instr_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_instr_MPORT_data = io_enq_bits_instr;
  assign ram_instr_MPORT_addr = enq_ptr_value;
  assign ram_instr_MPORT_mask = 1'h1;
  assign ram_instr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_pc_io_deq_bits_MPORT_en = 1'h1;
  assign ram_pc_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_pc_io_deq_bits_MPORT_data = ram_pc[ram_pc_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_pc_MPORT_data = io_enq_bits_pc;
  assign ram_pc_MPORT_addr = enq_ptr_value;
  assign ram_pc_MPORT_mask = 1'h1;
  assign ram_pc_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_pnpc_io_deq_bits_MPORT_en = 1'h1;
  assign ram_pnpc_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_pnpc_io_deq_bits_MPORT_data = ram_pnpc[ram_pnpc_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_pnpc_MPORT_data = io_enq_bits_pnpc;
  assign ram_pnpc_MPORT_addr = enq_ptr_value;
  assign ram_pnpc_MPORT_mask = 1'h1;
  assign ram_pnpc_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_0_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_0_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_0_io_deq_bits_MPORT_data = ram_exceptionVec_0[ram_exceptionVec_0_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_0_MPORT_data = 1'h0;
  assign ram_exceptionVec_0_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_0_MPORT_mask = 1'h1;
  assign ram_exceptionVec_0_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_1_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_1_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_1_io_deq_bits_MPORT_data = ram_exceptionVec_1[ram_exceptionVec_1_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_1_MPORT_data = io_enq_bits_exceptionVec_1;
  assign ram_exceptionVec_1_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_1_MPORT_mask = 1'h1;
  assign ram_exceptionVec_1_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_2_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_2_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_2_io_deq_bits_MPORT_data = ram_exceptionVec_2[ram_exceptionVec_2_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_2_MPORT_data = 1'h0;
  assign ram_exceptionVec_2_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_2_MPORT_mask = 1'h1;
  assign ram_exceptionVec_2_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_3_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_3_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_3_io_deq_bits_MPORT_data = ram_exceptionVec_3[ram_exceptionVec_3_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_3_MPORT_data = 1'h0;
  assign ram_exceptionVec_3_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_3_MPORT_mask = 1'h1;
  assign ram_exceptionVec_3_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_4_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_4_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_4_io_deq_bits_MPORT_data = ram_exceptionVec_4[ram_exceptionVec_4_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_4_MPORT_data = 1'h0;
  assign ram_exceptionVec_4_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_4_MPORT_mask = 1'h1;
  assign ram_exceptionVec_4_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_5_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_5_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_5_io_deq_bits_MPORT_data = ram_exceptionVec_5[ram_exceptionVec_5_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_5_MPORT_data = 1'h0;
  assign ram_exceptionVec_5_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_5_MPORT_mask = 1'h1;
  assign ram_exceptionVec_5_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_6_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_6_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_6_io_deq_bits_MPORT_data = ram_exceptionVec_6[ram_exceptionVec_6_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_6_MPORT_data = 1'h0;
  assign ram_exceptionVec_6_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_6_MPORT_mask = 1'h1;
  assign ram_exceptionVec_6_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_7_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_7_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_7_io_deq_bits_MPORT_data = ram_exceptionVec_7[ram_exceptionVec_7_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_7_MPORT_data = 1'h0;
  assign ram_exceptionVec_7_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_7_MPORT_mask = 1'h1;
  assign ram_exceptionVec_7_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_8_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_8_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_8_io_deq_bits_MPORT_data = ram_exceptionVec_8[ram_exceptionVec_8_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_8_MPORT_data = 1'h0;
  assign ram_exceptionVec_8_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_8_MPORT_mask = 1'h1;
  assign ram_exceptionVec_8_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_9_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_9_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_9_io_deq_bits_MPORT_data = ram_exceptionVec_9[ram_exceptionVec_9_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_9_MPORT_data = 1'h0;
  assign ram_exceptionVec_9_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_9_MPORT_mask = 1'h1;
  assign ram_exceptionVec_9_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_10_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_10_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_10_io_deq_bits_MPORT_data = ram_exceptionVec_10[ram_exceptionVec_10_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_10_MPORT_data = 1'h0;
  assign ram_exceptionVec_10_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_10_MPORT_mask = 1'h1;
  assign ram_exceptionVec_10_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_11_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_11_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_11_io_deq_bits_MPORT_data = ram_exceptionVec_11[ram_exceptionVec_11_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_11_MPORT_data = 1'h0;
  assign ram_exceptionVec_11_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_11_MPORT_mask = 1'h1;
  assign ram_exceptionVec_11_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_12_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_12_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_12_io_deq_bits_MPORT_data = ram_exceptionVec_12[ram_exceptionVec_12_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_12_MPORT_data = 1'h0;
  assign ram_exceptionVec_12_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_12_MPORT_mask = 1'h1;
  assign ram_exceptionVec_12_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_13_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_13_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_13_io_deq_bits_MPORT_data = ram_exceptionVec_13[ram_exceptionVec_13_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_13_MPORT_data = 1'h0;
  assign ram_exceptionVec_13_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_13_MPORT_mask = 1'h1;
  assign ram_exceptionVec_13_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_14_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_14_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_14_io_deq_bits_MPORT_data = ram_exceptionVec_14[ram_exceptionVec_14_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_14_MPORT_data = 1'h0;
  assign ram_exceptionVec_14_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_14_MPORT_mask = 1'h1;
  assign ram_exceptionVec_14_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_15_io_deq_bits_MPORT_en = 1'h1;
  assign ram_exceptionVec_15_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_exceptionVec_15_io_deq_bits_MPORT_data = ram_exceptionVec_15[ram_exceptionVec_15_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_exceptionVec_15_MPORT_data = 1'h0;
  assign ram_exceptionVec_15_MPORT_addr = enq_ptr_value;
  assign ram_exceptionVec_15_MPORT_mask = 1'h1;
  assign ram_exceptionVec_15_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_brIdx_io_deq_bits_MPORT_en = 1'h1;
  assign ram_brIdx_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_brIdx_io_deq_bits_MPORT_data = ram_brIdx[ram_brIdx_io_deq_bits_MPORT_addr]; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
  assign ram_brIdx_MPORT_data = io_enq_bits_brIdx;
  assign ram_brIdx_MPORT_addr = enq_ptr_value;
  assign ram_brIdx_MPORT_mask = 1'h1;
  assign ram_brIdx_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[src/main/scala/utils/FlushableQueue.scala 46:19]
  assign io_deq_valid = ~empty; // @[src/main/scala/utils/FlushableQueue.scala 45:19]
  assign io_deq_bits_instr = ram_instr_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_pc = ram_pc_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_pnpc = ram_pnpc_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_0 = ram_exceptionVec_0_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_1 = ram_exceptionVec_1_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_2 = ram_exceptionVec_2_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_3 = ram_exceptionVec_3_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_4 = ram_exceptionVec_4_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_5 = ram_exceptionVec_5_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_6 = ram_exceptionVec_6_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_7 = ram_exceptionVec_7_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_8 = ram_exceptionVec_8_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_9 = ram_exceptionVec_9_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_10 = ram_exceptionVec_10_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_11 = ram_exceptionVec_11_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_12 = ram_exceptionVec_12_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_13 = ram_exceptionVec_13_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_14 = ram_exceptionVec_14_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_exceptionVec_15 = ram_exceptionVec_15_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign io_deq_bits_brIdx = ram_brIdx_io_deq_bits_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 47:15]
  assign toggle_349_clock = clock;
  assign toggle_349_reset = reset;
  assign toggle_349_valid = enq_ptr_value ^ toggle_349_valid_reg;
  assign toggle_351_clock = clock;
  assign toggle_351_reset = reset;
  assign toggle_351_valid = deq_ptr_value ^ toggle_351_valid_reg;
  assign toggle_353_clock = clock;
  assign toggle_353_reset = reset;
  assign toggle_353_valid = maybe_full ^ toggle_353_valid_reg;
  always @(posedge clock) begin
    if (ram_instr_MPORT_en & ram_instr_MPORT_mask) begin
      ram_instr[ram_instr_MPORT_addr] <= ram_instr_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_pc_MPORT_en & ram_pc_MPORT_mask) begin
      ram_pc[ram_pc_MPORT_addr] <= ram_pc_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_pnpc_MPORT_en & ram_pnpc_MPORT_mask) begin
      ram_pnpc[ram_pnpc_MPORT_addr] <= ram_pnpc_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_0_MPORT_en & ram_exceptionVec_0_MPORT_mask) begin
      ram_exceptionVec_0[ram_exceptionVec_0_MPORT_addr] <= ram_exceptionVec_0_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_1_MPORT_en & ram_exceptionVec_1_MPORT_mask) begin
      ram_exceptionVec_1[ram_exceptionVec_1_MPORT_addr] <= ram_exceptionVec_1_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_2_MPORT_en & ram_exceptionVec_2_MPORT_mask) begin
      ram_exceptionVec_2[ram_exceptionVec_2_MPORT_addr] <= ram_exceptionVec_2_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_3_MPORT_en & ram_exceptionVec_3_MPORT_mask) begin
      ram_exceptionVec_3[ram_exceptionVec_3_MPORT_addr] <= ram_exceptionVec_3_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_4_MPORT_en & ram_exceptionVec_4_MPORT_mask) begin
      ram_exceptionVec_4[ram_exceptionVec_4_MPORT_addr] <= ram_exceptionVec_4_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_5_MPORT_en & ram_exceptionVec_5_MPORT_mask) begin
      ram_exceptionVec_5[ram_exceptionVec_5_MPORT_addr] <= ram_exceptionVec_5_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_6_MPORT_en & ram_exceptionVec_6_MPORT_mask) begin
      ram_exceptionVec_6[ram_exceptionVec_6_MPORT_addr] <= ram_exceptionVec_6_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_7_MPORT_en & ram_exceptionVec_7_MPORT_mask) begin
      ram_exceptionVec_7[ram_exceptionVec_7_MPORT_addr] <= ram_exceptionVec_7_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_8_MPORT_en & ram_exceptionVec_8_MPORT_mask) begin
      ram_exceptionVec_8[ram_exceptionVec_8_MPORT_addr] <= ram_exceptionVec_8_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_9_MPORT_en & ram_exceptionVec_9_MPORT_mask) begin
      ram_exceptionVec_9[ram_exceptionVec_9_MPORT_addr] <= ram_exceptionVec_9_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_10_MPORT_en & ram_exceptionVec_10_MPORT_mask) begin
      ram_exceptionVec_10[ram_exceptionVec_10_MPORT_addr] <= ram_exceptionVec_10_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_11_MPORT_en & ram_exceptionVec_11_MPORT_mask) begin
      ram_exceptionVec_11[ram_exceptionVec_11_MPORT_addr] <= ram_exceptionVec_11_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_12_MPORT_en & ram_exceptionVec_12_MPORT_mask) begin
      ram_exceptionVec_12[ram_exceptionVec_12_MPORT_addr] <= ram_exceptionVec_12_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_13_MPORT_en & ram_exceptionVec_13_MPORT_mask) begin
      ram_exceptionVec_13[ram_exceptionVec_13_MPORT_addr] <= ram_exceptionVec_13_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_14_MPORT_en & ram_exceptionVec_14_MPORT_mask) begin
      ram_exceptionVec_14[ram_exceptionVec_14_MPORT_addr] <= ram_exceptionVec_14_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_exceptionVec_15_MPORT_en & ram_exceptionVec_15_MPORT_mask) begin
      ram_exceptionVec_15[ram_exceptionVec_15_MPORT_addr] <= ram_exceptionVec_15_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (ram_brIdx_MPORT_en & ram_brIdx_MPORT_mask) begin
      ram_brIdx[ram_brIdx_MPORT_addr] <= ram_brIdx_MPORT_data; // @[src/main/scala/utils/FlushableQueue.scala 23:24]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (io_flush) begin // @[src/main/scala/utils/FlushableQueue.scala 62:19]
      enq_ptr_value <= 2'h0; // @[src/main/scala/utils/FlushableQueue.scala 64:21]
    end else if (do_enq) begin // @[src/main/scala/utils/FlushableQueue.scala 34:17]
      enq_ptr_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (io_flush) begin // @[src/main/scala/utils/FlushableQueue.scala 62:19]
      deq_ptr_value <= 2'h0; // @[src/main/scala/utils/FlushableQueue.scala 65:21]
    end else if (do_deq) begin // @[src/main/scala/utils/FlushableQueue.scala 38:17]
      deq_ptr_value <= _value_T_3; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/utils/FlushableQueue.scala 26:35]
      maybe_full <= 1'h0; // @[src/main/scala/utils/FlushableQueue.scala 26:35]
    end else if (io_flush) begin // @[src/main/scala/utils/FlushableQueue.scala 62:19]
      maybe_full <= 1'h0; // @[src/main/scala/utils/FlushableQueue.scala 67:16]
    end else if (do_enq != do_deq) begin // @[src/main/scala/utils/FlushableQueue.scala 41:28]
      maybe_full <= do_enq; // @[src/main/scala/utils/FlushableQueue.scala 42:16]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    enq_ptr_value_p <= enq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    toggle_349_valid_reg <= enq_ptr_value;
    deq_ptr_value_p <= deq_ptr_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    toggle_351_valid_reg <= deq_ptr_value;
    maybe_full_p <= maybe_full; // @[src/main/scala/utils/FlushableQueue.scala 26:35]
    toggle_353_valid_reg <= maybe_full;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_instr[initvar] = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_pc[initvar] = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_pnpc[initvar] = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_0[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_1[initvar] = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_2[initvar] = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_3[initvar] = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_4[initvar] = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_5[initvar] = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_6[initvar] = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_7[initvar] = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_8[initvar] = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_9[initvar] = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_10[initvar] = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_11[initvar] = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_12[initvar] = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_13[initvar] = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_14[initvar] = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_15[initvar] = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_brIdx[initvar] = _RAND_19[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  enq_ptr_value = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  deq_ptr_value = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  maybe_full = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  enq_ptr_value_p = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  toggle_349_valid_reg = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  deq_ptr_value_p = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  toggle_351_valid_reg = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  maybe_full_p = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  toggle_353_valid_reg = _RAND_28[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(enq_ptr_value_t[0]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(enq_ptr_value_t[1]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(deq_ptr_value_t[0]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(deq_ptr_value_t[1]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(maybe_full_t); // @[src/main/scala/utils/FlushableQueue.scala 26:35]
    end
  end
endmodule
module Frontend_inorder(
  input         clock,
  input         reset,
  input         io_imem_req_ready, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_imem_req_valid, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [38:0] io_imem_req_bits_addr, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [86:0] io_imem_req_bits_user, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_imem_resp_ready, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         io_imem_resp_valid, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input  [63:0] io_imem_resp_bits_rdata, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input  [86:0] io_imem_resp_bits_user, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         io_out_0_ready, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_valid, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [63:0] io_out_0_bits_cf_instr, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [38:0] io_out_0_bits_cf_pc, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [38:0] io_out_0_bits_cf_pnpc, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_intrVec_1, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_intrVec_3, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_intrVec_5, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_intrVec_7, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_intrVec_9, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_intrVec_11, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [3:0]  io_out_0_bits_cf_brIdx, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_ctrl_src1Type, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_ctrl_src2Type, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [2:0]  io_out_0_bits_ctrl_fuType, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [6:0]  io_out_0_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [4:0]  io_out_0_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [4:0]  io_out_0_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_ctrl_rfWen, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [4:0]  io_out_0_bits_ctrl_rfDest, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output        io_out_0_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [63:0] io_out_0_bits_data_imm, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  output [3:0]  io_flushVec, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input  [38:0] io_redirect_target, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         io_redirect_valid, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         io_iaf, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         io_sfence_vma_invalid, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         io_wfi_invalid, // @[src/main/scala/nutcore/frontend/Frontend.scala 41:14]
  input         REG_valid,
  input  [38:0] REG_pc,
  input         REG_isMissPredict,
  input  [38:0] REG_actualTarget,
  input  [6:0]  REG_fuOpType,
  input  [1:0]  REG_btbType,
  input         REG_isRVC,
  output        isWFI,
  input         flushICache,
  input         flushTLB,
  input  [11:0] intrVecIDU
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  wire  ifu_clock; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_reset; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_imem_req_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_imem_req_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [38:0] ifu_io_imem_req_bits_addr; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [81:0] ifu_io_imem_req_bits_user; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_imem_resp_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_imem_resp_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [63:0] ifu_io_imem_resp_bits_rdata; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [81:0] ifu_io_imem_resp_bits_user; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_out_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_out_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [63:0] ifu_io_out_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [38:0] ifu_io_out_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [38:0] ifu_io_out_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_out_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [3:0] ifu_io_out_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [38:0] ifu_io_redirect_target; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_redirect_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [3:0] ifu_io_flushVec; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_io_iaf; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_REG_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [38:0] ifu_REG_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_REG_isMissPredict; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [38:0] ifu_REG_actualTarget; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [6:0] ifu_REG_fuOpType; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire [1:0] ifu_REG_btbType; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_REG_isRVC; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_flushICache; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ifu_flushTLB; // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
  wire  ibf_clock; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_reset; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [63:0] ibf_io_in_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [38:0] ibf_io_in_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [38:0] ibf_io_in_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_0; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_3; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_4; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_6; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_8; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_9; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_10; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_13; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_14; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_in_bits_exceptionVec_15; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [3:0] ibf_io_in_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_out_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_out_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [63:0] ibf_io_out_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [38:0] ibf_io_out_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [38:0] ibf_io_out_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_out_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_out_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire [3:0] ibf_io_out_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_out_bits_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  ibf_io_flush; // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
  wire  idu_clock; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_reset; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_in_0_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_in_0_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [63:0] idu_io_in_0_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [38:0] idu_io_in_0_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [38:0] idu_io_in_0_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_in_0_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_in_0_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [3:0] idu_io_in_0_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_in_0_bits_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [63:0] idu_io_out_0_bits_cf_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [38:0] idu_io_out_0_bits_cf_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [38:0] idu_io_out_0_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [3:0] idu_io_out_0_bits_cf_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [2:0] idu_io_out_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [6:0] idu_io_out_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_out_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [63:0] idu_io_out_0_bits_data_imm; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_sfence_vma_invalid; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_io_wfi_invalid; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  idu_isWFI_0; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire [11:0] idu_intrVecIDU; // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
  wire  ibf_io_in_q_clock; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_reset; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_enq_ready; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_enq_valid; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [63:0] ibf_io_in_q_io_enq_bits_instr; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [38:0] ibf_io_in_q_io_enq_bits_pc; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [38:0] ibf_io_in_q_io_enq_bits_pnpc; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_enq_bits_exceptionVec_1; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [3:0] ibf_io_in_q_io_enq_bits_brIdx; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_ready; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_valid; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [63:0] ibf_io_in_q_io_deq_bits_instr; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [38:0] ibf_io_in_q_io_deq_bits_pc; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [38:0] ibf_io_in_q_io_deq_bits_pnpc; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_0; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_1; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_2; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_3; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_4; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_5; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_6; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_7; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_8; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_9; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_10; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_11; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_12; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_13; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_14; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_deq_bits_exceptionVec_15; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire [3:0] ibf_io_in_q_io_deq_bits_brIdx; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  ibf_io_in_q_io_flush; // @[src/main/scala/utils/FlushableQueue.scala 94:21]
  wire  _T_1 = idu_io_out_0_ready & idu_io_out_0_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  valid; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _GEN_0 = _T_1 ? 1'h0 : valid; // @[src/main/scala/utils/Pipeline.scala 24:24 25:{25,33}]
  wire  _T_3 = ibf_io_out_valid & idu_io_in_0_ready; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  _GEN_1 = ibf_io_out_valid & idu_io_in_0_ready | _GEN_0; // @[src/main/scala/utils/Pipeline.scala 26:{38,46}]
  reg [63:0] idu_io_in_0_bits_r_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] idu_io_in_0_bits_r_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] idu_io_in_0_bits_r_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  idu_io_in_0_bits_r_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  idu_io_in_0_bits_r_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] idu_io_in_0_bits_r_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  idu_io_in_0_bits_r_crossBoundaryFault; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  valid_p; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  valid_t = valid ^ valid_p; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  toggle_354_clock;
  wire  toggle_354_reset;
  wire  toggle_354_valid;
  reg  toggle_354_valid_reg;
  reg [63:0] idu_io_in_0_bits_r_instr_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [63:0] idu_io_in_0_bits_r_instr_t = idu_io_in_0_bits_r_instr ^ idu_io_in_0_bits_r_instr_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_355_clock;
  wire  toggle_355_reset;
  wire [63:0] toggle_355_valid;
  reg [63:0] toggle_355_valid_reg;
  reg [38:0] idu_io_in_0_bits_r_pc_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [38:0] idu_io_in_0_bits_r_pc_t = idu_io_in_0_bits_r_pc ^ idu_io_in_0_bits_r_pc_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_419_clock;
  wire  toggle_419_reset;
  wire [38:0] toggle_419_valid;
  reg [38:0] toggle_419_valid_reg;
  reg [38:0] idu_io_in_0_bits_r_pnpc_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [38:0] idu_io_in_0_bits_r_pnpc_t = idu_io_in_0_bits_r_pnpc ^ idu_io_in_0_bits_r_pnpc_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_458_clock;
  wire  toggle_458_reset;
  wire [38:0] toggle_458_valid;
  reg [38:0] toggle_458_valid_reg;
  reg  idu_io_in_0_bits_r_exceptionVec_1_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  idu_io_in_0_bits_r_exceptionVec_1_t = idu_io_in_0_bits_r_exceptionVec_1 ^ idu_io_in_0_bits_r_exceptionVec_1_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_497_clock;
  wire  toggle_497_reset;
  wire  toggle_497_valid;
  reg  toggle_497_valid_reg;
  reg  idu_io_in_0_bits_r_exceptionVec_12_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  idu_io_in_0_bits_r_exceptionVec_12_t = idu_io_in_0_bits_r_exceptionVec_12 ^ idu_io_in_0_bits_r_exceptionVec_12_p
    ; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_498_clock;
  wire  toggle_498_reset;
  wire  toggle_498_valid;
  reg  toggle_498_valid_reg;
  reg [3:0] idu_io_in_0_bits_r_brIdx_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [3:0] idu_io_in_0_bits_r_brIdx_t = idu_io_in_0_bits_r_brIdx ^ idu_io_in_0_bits_r_brIdx_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_499_clock;
  wire  toggle_499_reset;
  wire [3:0] toggle_499_valid;
  reg [3:0] toggle_499_valid_reg;
  reg  idu_io_in_0_bits_r_crossBoundaryFault_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  idu_io_in_0_bits_r_crossBoundaryFault_t = idu_io_in_0_bits_r_crossBoundaryFault ^
    idu_io_in_0_bits_r_crossBoundaryFault_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_503_clock;
  wire  toggle_503_reset;
  wire  toggle_503_valid;
  reg  toggle_503_valid_reg;
  IFU_inorder ifu ( // @[src/main/scala/nutcore/frontend/Frontend.scala 99:20]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_imem_req_ready(ifu_io_imem_req_ready),
    .io_imem_req_valid(ifu_io_imem_req_valid),
    .io_imem_req_bits_addr(ifu_io_imem_req_bits_addr),
    .io_imem_req_bits_user(ifu_io_imem_req_bits_user),
    .io_imem_resp_ready(ifu_io_imem_resp_ready),
    .io_imem_resp_valid(ifu_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(ifu_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(ifu_io_imem_resp_bits_user),
    .io_out_ready(ifu_io_out_ready),
    .io_out_valid(ifu_io_out_valid),
    .io_out_bits_instr(ifu_io_out_bits_instr),
    .io_out_bits_pc(ifu_io_out_bits_pc),
    .io_out_bits_pnpc(ifu_io_out_bits_pnpc),
    .io_out_bits_exceptionVec_1(ifu_io_out_bits_exceptionVec_1),
    .io_out_bits_brIdx(ifu_io_out_bits_brIdx),
    .io_redirect_target(ifu_io_redirect_target),
    .io_redirect_valid(ifu_io_redirect_valid),
    .io_flushVec(ifu_io_flushVec),
    .io_iaf(ifu_io_iaf),
    .REG_valid(ifu_REG_valid),
    .REG_pc(ifu_REG_pc),
    .REG_isMissPredict(ifu_REG_isMissPredict),
    .REG_actualTarget(ifu_REG_actualTarget),
    .REG_fuOpType(ifu_REG_fuOpType),
    .REG_btbType(ifu_REG_btbType),
    .REG_isRVC(ifu_REG_isRVC),
    .flushICache(ifu_flushICache),
    .flushTLB(ifu_flushTLB)
  );
  NaiveRVCAlignBuffer ibf ( // @[src/main/scala/nutcore/frontend/Frontend.scala 100:19]
    .clock(ibf_clock),
    .reset(ibf_reset),
    .io_in_ready(ibf_io_in_ready),
    .io_in_valid(ibf_io_in_valid),
    .io_in_bits_instr(ibf_io_in_bits_instr),
    .io_in_bits_pc(ibf_io_in_bits_pc),
    .io_in_bits_pnpc(ibf_io_in_bits_pnpc),
    .io_in_bits_exceptionVec_0(ibf_io_in_bits_exceptionVec_0),
    .io_in_bits_exceptionVec_1(ibf_io_in_bits_exceptionVec_1),
    .io_in_bits_exceptionVec_2(ibf_io_in_bits_exceptionVec_2),
    .io_in_bits_exceptionVec_3(ibf_io_in_bits_exceptionVec_3),
    .io_in_bits_exceptionVec_4(ibf_io_in_bits_exceptionVec_4),
    .io_in_bits_exceptionVec_5(ibf_io_in_bits_exceptionVec_5),
    .io_in_bits_exceptionVec_6(ibf_io_in_bits_exceptionVec_6),
    .io_in_bits_exceptionVec_7(ibf_io_in_bits_exceptionVec_7),
    .io_in_bits_exceptionVec_8(ibf_io_in_bits_exceptionVec_8),
    .io_in_bits_exceptionVec_9(ibf_io_in_bits_exceptionVec_9),
    .io_in_bits_exceptionVec_10(ibf_io_in_bits_exceptionVec_10),
    .io_in_bits_exceptionVec_11(ibf_io_in_bits_exceptionVec_11),
    .io_in_bits_exceptionVec_12(ibf_io_in_bits_exceptionVec_12),
    .io_in_bits_exceptionVec_13(ibf_io_in_bits_exceptionVec_13),
    .io_in_bits_exceptionVec_14(ibf_io_in_bits_exceptionVec_14),
    .io_in_bits_exceptionVec_15(ibf_io_in_bits_exceptionVec_15),
    .io_in_bits_brIdx(ibf_io_in_bits_brIdx),
    .io_out_ready(ibf_io_out_ready),
    .io_out_valid(ibf_io_out_valid),
    .io_out_bits_instr(ibf_io_out_bits_instr),
    .io_out_bits_pc(ibf_io_out_bits_pc),
    .io_out_bits_pnpc(ibf_io_out_bits_pnpc),
    .io_out_bits_exceptionVec_1(ibf_io_out_bits_exceptionVec_1),
    .io_out_bits_exceptionVec_12(ibf_io_out_bits_exceptionVec_12),
    .io_out_bits_brIdx(ibf_io_out_bits_brIdx),
    .io_out_bits_crossBoundaryFault(ibf_io_out_bits_crossBoundaryFault),
    .io_flush(ibf_io_flush)
  );
  IDU idu ( // @[src/main/scala/nutcore/frontend/Frontend.scala 101:20]
    .clock(idu_clock),
    .reset(idu_reset),
    .io_in_0_ready(idu_io_in_0_ready),
    .io_in_0_valid(idu_io_in_0_valid),
    .io_in_0_bits_instr(idu_io_in_0_bits_instr),
    .io_in_0_bits_pc(idu_io_in_0_bits_pc),
    .io_in_0_bits_pnpc(idu_io_in_0_bits_pnpc),
    .io_in_0_bits_exceptionVec_1(idu_io_in_0_bits_exceptionVec_1),
    .io_in_0_bits_exceptionVec_12(idu_io_in_0_bits_exceptionVec_12),
    .io_in_0_bits_brIdx(idu_io_in_0_bits_brIdx),
    .io_in_0_bits_crossBoundaryFault(idu_io_in_0_bits_crossBoundaryFault),
    .io_out_0_ready(idu_io_out_0_ready),
    .io_out_0_valid(idu_io_out_0_valid),
    .io_out_0_bits_cf_instr(idu_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(idu_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(idu_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(idu_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(idu_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(idu_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_intrVec_1(idu_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_3(idu_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_5(idu_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_7(idu_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_9(idu_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_11(idu_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(idu_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_cf_crossBoundaryFault(idu_io_out_0_bits_cf_crossBoundaryFault),
    .io_out_0_bits_ctrl_src1Type(idu_io_out_0_bits_ctrl_src1Type),
    .io_out_0_bits_ctrl_src2Type(idu_io_out_0_bits_ctrl_src2Type),
    .io_out_0_bits_ctrl_fuType(idu_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(idu_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfSrc1(idu_io_out_0_bits_ctrl_rfSrc1),
    .io_out_0_bits_ctrl_rfSrc2(idu_io_out_0_bits_ctrl_rfSrc2),
    .io_out_0_bits_ctrl_rfWen(idu_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(idu_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_ctrl_isNutCoreTrap(idu_io_out_0_bits_ctrl_isNutCoreTrap),
    .io_out_0_bits_data_imm(idu_io_out_0_bits_data_imm),
    .io_sfence_vma_invalid(idu_io_sfence_vma_invalid),
    .io_wfi_invalid(idu_io_wfi_invalid),
    .isWFI_0(idu_isWFI_0),
    .intrVecIDU(idu_intrVecIDU)
  );
  FlushableQueue ibf_io_in_q ( // @[src/main/scala/utils/FlushableQueue.scala 94:21]
    .clock(ibf_io_in_q_clock),
    .reset(ibf_io_in_q_reset),
    .io_enq_ready(ibf_io_in_q_io_enq_ready),
    .io_enq_valid(ibf_io_in_q_io_enq_valid),
    .io_enq_bits_instr(ibf_io_in_q_io_enq_bits_instr),
    .io_enq_bits_pc(ibf_io_in_q_io_enq_bits_pc),
    .io_enq_bits_pnpc(ibf_io_in_q_io_enq_bits_pnpc),
    .io_enq_bits_exceptionVec_1(ibf_io_in_q_io_enq_bits_exceptionVec_1),
    .io_enq_bits_brIdx(ibf_io_in_q_io_enq_bits_brIdx),
    .io_deq_ready(ibf_io_in_q_io_deq_ready),
    .io_deq_valid(ibf_io_in_q_io_deq_valid),
    .io_deq_bits_instr(ibf_io_in_q_io_deq_bits_instr),
    .io_deq_bits_pc(ibf_io_in_q_io_deq_bits_pc),
    .io_deq_bits_pnpc(ibf_io_in_q_io_deq_bits_pnpc),
    .io_deq_bits_exceptionVec_0(ibf_io_in_q_io_deq_bits_exceptionVec_0),
    .io_deq_bits_exceptionVec_1(ibf_io_in_q_io_deq_bits_exceptionVec_1),
    .io_deq_bits_exceptionVec_2(ibf_io_in_q_io_deq_bits_exceptionVec_2),
    .io_deq_bits_exceptionVec_3(ibf_io_in_q_io_deq_bits_exceptionVec_3),
    .io_deq_bits_exceptionVec_4(ibf_io_in_q_io_deq_bits_exceptionVec_4),
    .io_deq_bits_exceptionVec_5(ibf_io_in_q_io_deq_bits_exceptionVec_5),
    .io_deq_bits_exceptionVec_6(ibf_io_in_q_io_deq_bits_exceptionVec_6),
    .io_deq_bits_exceptionVec_7(ibf_io_in_q_io_deq_bits_exceptionVec_7),
    .io_deq_bits_exceptionVec_8(ibf_io_in_q_io_deq_bits_exceptionVec_8),
    .io_deq_bits_exceptionVec_9(ibf_io_in_q_io_deq_bits_exceptionVec_9),
    .io_deq_bits_exceptionVec_10(ibf_io_in_q_io_deq_bits_exceptionVec_10),
    .io_deq_bits_exceptionVec_11(ibf_io_in_q_io_deq_bits_exceptionVec_11),
    .io_deq_bits_exceptionVec_12(ibf_io_in_q_io_deq_bits_exceptionVec_12),
    .io_deq_bits_exceptionVec_13(ibf_io_in_q_io_deq_bits_exceptionVec_13),
    .io_deq_bits_exceptionVec_14(ibf_io_in_q_io_deq_bits_exceptionVec_14),
    .io_deq_bits_exceptionVec_15(ibf_io_in_q_io_deq_bits_exceptionVec_15),
    .io_deq_bits_brIdx(ibf_io_in_q_io_deq_bits_brIdx),
    .io_flush(ibf_io_in_q_io_flush)
  );
  GEN_w1_toggle #(.COVER_INDEX(354)) toggle_354 (
    .clock(toggle_354_clock),
    .reset(toggle_354_reset),
    .valid(toggle_354_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(355)) toggle_355 (
    .clock(toggle_355_clock),
    .reset(toggle_355_reset),
    .valid(toggle_355_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(419)) toggle_419 (
    .clock(toggle_419_clock),
    .reset(toggle_419_reset),
    .valid(toggle_419_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(458)) toggle_458 (
    .clock(toggle_458_clock),
    .reset(toggle_458_reset),
    .valid(toggle_458_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(497)) toggle_497 (
    .clock(toggle_497_clock),
    .reset(toggle_497_reset),
    .valid(toggle_497_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(498)) toggle_498 (
    .clock(toggle_498_clock),
    .reset(toggle_498_reset),
    .valid(toggle_498_valid)
  );
  GEN_w4_toggle #(.COVER_INDEX(499)) toggle_499 (
    .clock(toggle_499_clock),
    .reset(toggle_499_reset),
    .valid(toggle_499_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(503)) toggle_503 (
    .clock(toggle_503_clock),
    .reset(toggle_503_reset),
    .valid(toggle_503_valid)
  );
  assign io_imem_req_valid = ifu_io_imem_req_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign io_imem_req_bits_addr = ifu_io_imem_req_bits_addr; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign io_imem_req_bits_user = {{5'd0}, ifu_io_imem_req_bits_user}; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign io_imem_resp_ready = ifu_io_imem_resp_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign io_out_0_valid = idu_io_out_0_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_instr = idu_io_out_0_bits_cf_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_pc = idu_io_out_0_bits_cf_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_pnpc = idu_io_out_0_bits_cf_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_exceptionVec_1 = idu_io_out_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_exceptionVec_2 = idu_io_out_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_exceptionVec_12 = idu_io_out_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_intrVec_1 = idu_io_out_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_intrVec_3 = idu_io_out_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_intrVec_5 = idu_io_out_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_intrVec_7 = idu_io_out_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_intrVec_9 = idu_io_out_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_intrVec_11 = idu_io_out_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_brIdx = idu_io_out_0_bits_cf_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_cf_crossBoundaryFault = idu_io_out_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_src1Type = idu_io_out_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_src2Type = idu_io_out_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_fuType = idu_io_out_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_fuOpType = idu_io_out_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_rfSrc1 = idu_io_out_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_rfSrc2 = idu_io_out_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_rfWen = idu_io_out_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_rfDest = idu_io_out_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_ctrl_isNutCoreTrap = idu_io_out_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_out_0_bits_data_imm = idu_io_out_0_bits_data_imm; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign io_flushVec = ifu_io_flushVec; // @[src/main/scala/nutcore/frontend/Frontend.scala 119:15]
  assign isWFI = idu_isWFI_0;
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_imem_req_ready = io_imem_req_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign ifu_io_imem_resp_valid = io_imem_resp_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign ifu_io_imem_resp_bits_rdata = io_imem_resp_bits_rdata; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign ifu_io_imem_resp_bits_user = io_imem_resp_bits_user[81:0]; // @[src/main/scala/nutcore/frontend/Frontend.scala 123:11]
  assign ifu_io_out_ready = ibf_io_in_q_io_enq_ready; // @[src/main/scala/utils/FlushableQueue.scala 98:17]
  assign ifu_io_redirect_target = io_redirect_target; // @[src/main/scala/nutcore/frontend/Frontend.scala 118:15]
  assign ifu_io_redirect_valid = io_redirect_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 118:15]
  assign ifu_io_iaf = io_iaf; // @[src/main/scala/nutcore/frontend/Frontend.scala 122:10]
  assign ifu_REG_valid = REG_valid;
  assign ifu_REG_pc = REG_pc;
  assign ifu_REG_isMissPredict = REG_isMissPredict;
  assign ifu_REG_actualTarget = REG_actualTarget;
  assign ifu_REG_fuOpType = REG_fuOpType;
  assign ifu_REG_btbType = REG_btbType;
  assign ifu_REG_isRVC = REG_isRVC;
  assign ifu_flushICache = flushICache;
  assign ifu_flushTLB = flushTLB;
  assign ibf_clock = clock;
  assign ibf_reset = reset;
  assign ibf_io_in_valid = ibf_io_in_q_io_deq_valid; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_instr = ibf_io_in_q_io_deq_bits_instr; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_pc = ibf_io_in_q_io_deq_bits_pc; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_pnpc = ibf_io_in_q_io_deq_bits_pnpc; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_0 = ibf_io_in_q_io_deq_bits_exceptionVec_0; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_1 = ibf_io_in_q_io_deq_bits_exceptionVec_1; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_2 = ibf_io_in_q_io_deq_bits_exceptionVec_2; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_3 = ibf_io_in_q_io_deq_bits_exceptionVec_3; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_4 = ibf_io_in_q_io_deq_bits_exceptionVec_4; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_5 = ibf_io_in_q_io_deq_bits_exceptionVec_5; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_6 = ibf_io_in_q_io_deq_bits_exceptionVec_6; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_7 = ibf_io_in_q_io_deq_bits_exceptionVec_7; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_8 = ibf_io_in_q_io_deq_bits_exceptionVec_8; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_9 = ibf_io_in_q_io_deq_bits_exceptionVec_9; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_10 = ibf_io_in_q_io_deq_bits_exceptionVec_10; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_11 = ibf_io_in_q_io_deq_bits_exceptionVec_11; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_12 = ibf_io_in_q_io_deq_bits_exceptionVec_12; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_13 = ibf_io_in_q_io_deq_bits_exceptionVec_13; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_14 = ibf_io_in_q_io_deq_bits_exceptionVec_14; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_exceptionVec_15 = ibf_io_in_q_io_deq_bits_exceptionVec_15; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_bits_brIdx = ibf_io_in_q_io_deq_bits_brIdx; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_out_ready = idu_io_in_0_ready; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign ibf_io_flush = ifu_io_flushVec[1]; // @[src/main/scala/nutcore/frontend/Frontend.scala 116:34]
  assign idu_clock = clock;
  assign idu_reset = reset;
  assign idu_io_in_0_valid = valid; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign idu_io_in_0_bits_instr = idu_io_in_0_bits_r_instr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_pc = idu_io_in_0_bits_r_pc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_pnpc = idu_io_in_0_bits_r_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_exceptionVec_1 = idu_io_in_0_bits_r_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_exceptionVec_12 = idu_io_in_0_bits_r_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_brIdx = idu_io_in_0_bits_r_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_in_0_bits_crossBoundaryFault = idu_io_in_0_bits_r_crossBoundaryFault; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign idu_io_out_0_ready = io_out_0_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 117:10]
  assign idu_io_sfence_vma_invalid = io_sfence_vma_invalid; // @[src/main/scala/nutcore/frontend/Frontend.scala 113:29]
  assign idu_io_wfi_invalid = io_wfi_invalid; // @[src/main/scala/nutcore/frontend/Frontend.scala 114:22]
  assign idu_intrVecIDU = intrVecIDU;
  assign ibf_io_in_q_clock = clock;
  assign ibf_io_in_q_reset = reset;
  assign ibf_io_in_q_io_enq_valid = ifu_io_out_valid; // @[src/main/scala/utils/FlushableQueue.scala 95:22]
  assign ibf_io_in_q_io_enq_bits_instr = ifu_io_out_bits_instr; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_enq_bits_pc = ifu_io_out_bits_pc; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_enq_bits_pnpc = ifu_io_out_bits_pnpc; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_enq_bits_exceptionVec_1 = ifu_io_out_bits_exceptionVec_1; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_enq_bits_brIdx = ifu_io_out_bits_brIdx; // @[src/main/scala/utils/FlushableQueue.scala 96:21]
  assign ibf_io_in_q_io_deq_ready = ibf_io_in_ready; // @[src/main/scala/nutcore/frontend/Frontend.scala 107:11]
  assign ibf_io_in_q_io_flush = ifu_io_flushVec[0]; // @[src/main/scala/nutcore/frontend/Frontend.scala 110:58]
  assign toggle_354_clock = clock;
  assign toggle_354_reset = reset;
  assign toggle_354_valid = valid ^ toggle_354_valid_reg;
  assign toggle_355_clock = clock;
  assign toggle_355_reset = reset;
  assign toggle_355_valid = idu_io_in_0_bits_r_instr ^ toggle_355_valid_reg;
  assign toggle_419_clock = clock;
  assign toggle_419_reset = reset;
  assign toggle_419_valid = idu_io_in_0_bits_r_pc ^ toggle_419_valid_reg;
  assign toggle_458_clock = clock;
  assign toggle_458_reset = reset;
  assign toggle_458_valid = idu_io_in_0_bits_r_pnpc ^ toggle_458_valid_reg;
  assign toggle_497_clock = clock;
  assign toggle_497_reset = reset;
  assign toggle_497_valid = idu_io_in_0_bits_r_exceptionVec_1 ^ toggle_497_valid_reg;
  assign toggle_498_clock = clock;
  assign toggle_498_reset = reset;
  assign toggle_498_valid = idu_io_in_0_bits_r_exceptionVec_12 ^ toggle_498_valid_reg;
  assign toggle_499_clock = clock;
  assign toggle_499_reset = reset;
  assign toggle_499_valid = idu_io_in_0_bits_r_brIdx ^ toggle_499_valid_reg;
  assign toggle_503_clock = clock;
  assign toggle_503_reset = reset;
  assign toggle_503_valid = idu_io_in_0_bits_r_crossBoundaryFault ^ toggle_503_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else if (ifu_io_flushVec[1]) begin // @[src/main/scala/utils/Pipeline.scala 27:20]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 27:28]
    end else begin
      valid <= _GEN_1;
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_instr <= ibf_io_out_bits_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_pc <= ibf_io_out_bits_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_pnpc <= ibf_io_out_bits_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_exceptionVec_1 <= ibf_io_out_bits_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_exceptionVec_12 <= ibf_io_out_bits_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_brIdx <= ibf_io_out_bits_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_3) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      idu_io_in_0_bits_r_crossBoundaryFault <= ibf_io_out_bits_crossBoundaryFault; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    valid_p <= valid; // @[src/main/scala/utils/Pipeline.scala 24:24]
    toggle_354_valid_reg <= valid;
    idu_io_in_0_bits_r_instr_p <= idu_io_in_0_bits_r_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_355_valid_reg <= idu_io_in_0_bits_r_instr;
    idu_io_in_0_bits_r_pc_p <= idu_io_in_0_bits_r_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_419_valid_reg <= idu_io_in_0_bits_r_pc;
    idu_io_in_0_bits_r_pnpc_p <= idu_io_in_0_bits_r_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_458_valid_reg <= idu_io_in_0_bits_r_pnpc;
    idu_io_in_0_bits_r_exceptionVec_1_p <= idu_io_in_0_bits_r_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_497_valid_reg <= idu_io_in_0_bits_r_exceptionVec_1;
    idu_io_in_0_bits_r_exceptionVec_12_p <= idu_io_in_0_bits_r_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_498_valid_reg <= idu_io_in_0_bits_r_exceptionVec_12;
    idu_io_in_0_bits_r_brIdx_p <= idu_io_in_0_bits_r_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_499_valid_reg <= idu_io_in_0_bits_r_brIdx;
    idu_io_in_0_bits_r_crossBoundaryFault_p <= idu_io_in_0_bits_r_crossBoundaryFault; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_503_valid_reg <= idu_io_in_0_bits_r_crossBoundaryFault;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  idu_io_in_0_bits_r_instr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  idu_io_in_0_bits_r_pc = _RAND_2[38:0];
  _RAND_3 = {2{`RANDOM}};
  idu_io_in_0_bits_r_pnpc = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  idu_io_in_0_bits_r_exceptionVec_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  idu_io_in_0_bits_r_exceptionVec_12 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  idu_io_in_0_bits_r_brIdx = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  idu_io_in_0_bits_r_crossBoundaryFault = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  valid_p = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  toggle_354_valid_reg = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  idu_io_in_0_bits_r_instr_p = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  toggle_355_valid_reg = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  idu_io_in_0_bits_r_pc_p = _RAND_12[38:0];
  _RAND_13 = {2{`RANDOM}};
  toggle_419_valid_reg = _RAND_13[38:0];
  _RAND_14 = {2{`RANDOM}};
  idu_io_in_0_bits_r_pnpc_p = _RAND_14[38:0];
  _RAND_15 = {2{`RANDOM}};
  toggle_458_valid_reg = _RAND_15[38:0];
  _RAND_16 = {1{`RANDOM}};
  idu_io_in_0_bits_r_exceptionVec_1_p = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  toggle_497_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  idu_io_in_0_bits_r_exceptionVec_12_p = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  toggle_498_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  idu_io_in_0_bits_r_brIdx_p = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  toggle_499_valid_reg = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  idu_io_in_0_bits_r_crossBoundaryFault_p = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  toggle_503_valid_reg = _RAND_23[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(valid_t); // @[src/main/scala/utils/Pipeline.scala 24:24]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[5]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[6]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[7]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[8]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[9]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[10]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[11]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[12]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[13]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[14]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[15]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[16]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[17]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[18]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[19]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[20]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[21]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[22]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[23]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[24]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[25]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[26]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[27]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[28]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[29]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[30]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[31]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[32]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[33]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[34]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[35]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[36]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[37]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[38]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[39]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[40]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[41]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[42]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[43]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[44]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[45]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[46]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[47]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[48]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[49]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[50]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[51]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[52]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[53]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[54]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[55]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[56]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[57]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[58]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[59]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[60]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[61]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[62]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_instr_t[63]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[5]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[6]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[7]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[8]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[9]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[10]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[11]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[12]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[13]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[14]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[15]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[16]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[17]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[18]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[19]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[20]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[21]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[22]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[23]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[24]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[25]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[26]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[27]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[28]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[29]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[30]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[31]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[32]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[33]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[34]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[35]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[36]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[37]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pc_t[38]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[5]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[6]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[7]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[8]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[9]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[10]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[11]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[12]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[13]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[14]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[15]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[16]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[17]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[18]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[19]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[20]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[21]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[22]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[23]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[24]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[25]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[26]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[27]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[28]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[29]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[30]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[31]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[32]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[33]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[34]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[35]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[36]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[37]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_pnpc_t[38]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_exceptionVec_1_t); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_exceptionVec_12_t); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_brIdx_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_brIdx_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_brIdx_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_brIdx_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(idu_io_in_0_bits_r_crossBoundaryFault_t); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
  end
endmodule
module DummyDPICWrapper(
  input         clock,
  input         reset,
  input  [63:0] io_bits_value_1, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_2, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_3, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_4, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_5, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_6, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_7, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_8, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_9, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_10, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_11, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_12, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_13, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_14, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_15, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_16, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_17, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_18, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_19, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_20, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_21, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_22, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_23, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_24, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_25, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_26, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_27, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_28, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_29, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_30, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_value_31 // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_0; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_1; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_2; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_3; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_4; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_5; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_6; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_7; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_8; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_9; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_10; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_11; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_12; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_13; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_14; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_15; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_16; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_17; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_18; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_19; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_20; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_21; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_22; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_23; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_24; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_25; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_26; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_27; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_28; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_29; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_30; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_value_31; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestArchIntRegState dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_value_0(dpic_io_value_0),
    .io_value_1(dpic_io_value_1),
    .io_value_2(dpic_io_value_2),
    .io_value_3(dpic_io_value_3),
    .io_value_4(dpic_io_value_4),
    .io_value_5(dpic_io_value_5),
    .io_value_6(dpic_io_value_6),
    .io_value_7(dpic_io_value_7),
    .io_value_8(dpic_io_value_8),
    .io_value_9(dpic_io_value_9),
    .io_value_10(dpic_io_value_10),
    .io_value_11(dpic_io_value_11),
    .io_value_12(dpic_io_value_12),
    .io_value_13(dpic_io_value_13),
    .io_value_14(dpic_io_value_14),
    .io_value_15(dpic_io_value_15),
    .io_value_16(dpic_io_value_16),
    .io_value_17(dpic_io_value_17),
    .io_value_18(dpic_io_value_18),
    .io_value_19(dpic_io_value_19),
    .io_value_20(dpic_io_value_20),
    .io_value_21(dpic_io_value_21),
    .io_value_22(dpic_io_value_22),
    .io_value_23(dpic_io_value_23),
    .io_value_24(dpic_io_value_24),
    .io_value_25(dpic_io_value_25),
    .io_value_26(dpic_io_value_26),
    .io_value_27(dpic_io_value_27),
    .io_value_28(dpic_io_value_28),
    .io_value_29(dpic_io_value_29),
    .io_value_30(dpic_io_value_30),
    .io_value_31(dpic_io_value_31),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = 1'h1; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_value_0 = 64'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_1 = io_bits_value_1; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_2 = io_bits_value_2; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_3 = io_bits_value_3; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_4 = io_bits_value_4; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_5 = io_bits_value_5; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_6 = io_bits_value_6; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_7 = io_bits_value_7; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_8 = io_bits_value_8; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_9 = io_bits_value_9; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_10 = io_bits_value_10; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_11 = io_bits_value_11; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_12 = io_bits_value_12; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_13 = io_bits_value_13; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_14 = io_bits_value_14; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_15 = io_bits_value_15; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_16 = io_bits_value_16; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_17 = io_bits_value_17; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_18 = io_bits_value_18; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_19 = io_bits_value_19; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_20 = io_bits_value_20; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_21 = io_bits_value_21; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_22 = io_bits_value_22; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_23 = io_bits_value_23; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_24 = io_bits_value_24; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_25 = io_bits_value_25; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_26 = io_bits_value_26; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_27 = io_bits_value_27; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_28 = io_bits_value_28; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_29 = io_bits_value_29; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_30 = io_bits_value_30; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_value_31 = io_bits_value_31; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module ISU(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_valid, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [63:0] io_in_0_bits_cf_instr, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [38:0] io_in_0_bits_cf_pc, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [38:0] io_in_0_bits_cf_pnpc, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_3, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_5, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_7, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_9, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_intrVec_11, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [3:0]  io_in_0_bits_cf_brIdx, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_ctrl_src1Type, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_ctrl_src2Type, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [2:0]  io_in_0_bits_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [6:0]  io_in_0_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_in_0_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_in_0_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_in_0_bits_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_in_0_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [63:0] io_in_0_bits_data_imm, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [63:0] io_out_bits_cf_instr, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [38:0] io_out_bits_cf_pc, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [38:0] io_out_bits_cf_pnpc, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_3, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_5, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_7, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_9, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_intrVec_11, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [3:0]  io_out_bits_cf_brIdx, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [2:0]  io_out_bits_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [6:0]  io_out_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [4:0]  io_out_bits_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output        io_out_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [63:0] io_out_bits_data_src1, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [63:0] io_out_bits_data_src2, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  output [63:0] io_out_bits_data_imm, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_wb_rfWen, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_wb_rfDest, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [63:0] io_wb_rfData, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_forward_valid, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_forward_wb_rfWen, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [4:0]  io_forward_wb_rfDest, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [63:0] io_forward_wb_rfData, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input  [2:0]  io_forward_fuType, // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
  input         io_flush // @[src/main/scala/nutcore/backend/seq/ISU.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
`endif // RANDOMIZE_REG_INIT
  wire  difftest_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_1; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_2; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_3; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_4; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_5; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_6; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_7; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_8; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_9; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_10; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_11; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_12; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_13; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_14; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_15; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_16; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_17; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_18; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_19; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_20; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_21; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_22; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_23; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_24; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_25; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_26; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_27; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_28; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_29; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_30; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_value_31; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  forwardRfWen = io_forward_wb_rfWen & io_forward_valid; // @[src/main/scala/nutcore/backend/seq/ISU.scala 43:42]
  wire  dontForward1 = io_forward_fuType != 3'h0 & io_forward_fuType != 3'h1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 44:57]
  wire  src1DependEX = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_forward_wb_rfDest &
    forwardRfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire  src2DependEX = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_forward_wb_rfDest &
    forwardRfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire  src1DependWB = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_wb_rfDest & io_wb_rfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire  src2DependWB = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_wb_rfDest & io_wb_rfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire  _src1ForwardNextCycle_T = ~dontForward1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 50:46]
  wire  src1ForwardNextCycle = src1DependEX & ~dontForward1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 50:43]
  wire  src2ForwardNextCycle = src2DependEX & _src1ForwardNextCycle_T; // @[src/main/scala/nutcore/backend/seq/ISU.scala 51:43]
  wire  _src1Forward_T_1 = dontForward1 ? ~src1DependEX : 1'h1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 52:40]
  wire  src1Forward = src1DependWB & _src1Forward_T_1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 52:34]
  wire  _src2Forward_T_1 = dontForward1 ? ~src2DependEX : 1'h1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 53:40]
  wire  src2Forward = src2DependWB & _src2Forward_T_1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 53:34]
  reg [31:0] busy; // @[src/main/scala/nutcore/RF.scala 37:21]
  wire [31:0] _src1Ready_T = busy >> io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/RF.scala 38:37]
  wire  src1Ready = ~_src1Ready_T[0] | src1ForwardNextCycle | src1Forward; // @[src/main/scala/nutcore/backend/seq/ISU.scala 56:62]
  wire [31:0] _src2Ready_T = busy >> io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/RF.scala 38:37]
  wire  src2Ready = ~_src2Ready_T[0] | src2ForwardNextCycle | src2Forward; // @[src/main/scala/nutcore/backend/seq/ISU.scala 57:62]
  reg [63:0] rf_0; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_1; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_2; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_3; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_4; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_5; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_6; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_7; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_8; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_9; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_10; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_11; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_12; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_13; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_14; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_15; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_16; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_17; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_18; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_19; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_20; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_21; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_22; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_23; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_24; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_25; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_26; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_27; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_28; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_29; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_30; // @[src/main/scala/nutcore/RF.scala 31:19]
  reg [63:0] rf_31; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  io_out_bits_data_src1_signBit = io_in_0_bits_cf_pc[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _io_out_bits_data_src1_T_1 = io_out_bits_data_src1_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _io_out_bits_data_src1_T_2 = {_io_out_bits_data_src1_T_1,io_in_0_bits_cf_pc}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  _io_out_bits_data_src1_T_3 = ~src1ForwardNextCycle; // @[src/main/scala/nutcore/backend/seq/ISU.scala 66:21]
  wire  _io_out_bits_data_src1_T_4 = src1Forward & ~src1ForwardNextCycle; // @[src/main/scala/nutcore/backend/seq/ISU.scala 66:18]
  wire  _io_out_bits_data_src1_T_9 = ~io_in_0_bits_ctrl_src1Type & _io_out_bits_data_src1_T_3 & ~src1Forward; // @[src/main/scala/nutcore/backend/seq/ISU.scala 67:76]
  wire [63:0] _GEN_1 = 5'h1 == io_in_0_bits_ctrl_rfSrc1 ? rf_1 : rf_0; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_2 = 5'h2 == io_in_0_bits_ctrl_rfSrc1 ? rf_2 : _GEN_1; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_3 = 5'h3 == io_in_0_bits_ctrl_rfSrc1 ? rf_3 : _GEN_2; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_4 = 5'h4 == io_in_0_bits_ctrl_rfSrc1 ? rf_4 : _GEN_3; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_5 = 5'h5 == io_in_0_bits_ctrl_rfSrc1 ? rf_5 : _GEN_4; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_6 = 5'h6 == io_in_0_bits_ctrl_rfSrc1 ? rf_6 : _GEN_5; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_7 = 5'h7 == io_in_0_bits_ctrl_rfSrc1 ? rf_7 : _GEN_6; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_8 = 5'h8 == io_in_0_bits_ctrl_rfSrc1 ? rf_8 : _GEN_7; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_9 = 5'h9 == io_in_0_bits_ctrl_rfSrc1 ? rf_9 : _GEN_8; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_10 = 5'ha == io_in_0_bits_ctrl_rfSrc1 ? rf_10 : _GEN_9; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_11 = 5'hb == io_in_0_bits_ctrl_rfSrc1 ? rf_11 : _GEN_10; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_12 = 5'hc == io_in_0_bits_ctrl_rfSrc1 ? rf_12 : _GEN_11; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_13 = 5'hd == io_in_0_bits_ctrl_rfSrc1 ? rf_13 : _GEN_12; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_14 = 5'he == io_in_0_bits_ctrl_rfSrc1 ? rf_14 : _GEN_13; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_15 = 5'hf == io_in_0_bits_ctrl_rfSrc1 ? rf_15 : _GEN_14; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_16 = 5'h10 == io_in_0_bits_ctrl_rfSrc1 ? rf_16 : _GEN_15; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_17 = 5'h11 == io_in_0_bits_ctrl_rfSrc1 ? rf_17 : _GEN_16; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_18 = 5'h12 == io_in_0_bits_ctrl_rfSrc1 ? rf_18 : _GEN_17; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_19 = 5'h13 == io_in_0_bits_ctrl_rfSrc1 ? rf_19 : _GEN_18; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_20 = 5'h14 == io_in_0_bits_ctrl_rfSrc1 ? rf_20 : _GEN_19; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_21 = 5'h15 == io_in_0_bits_ctrl_rfSrc1 ? rf_21 : _GEN_20; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_22 = 5'h16 == io_in_0_bits_ctrl_rfSrc1 ? rf_22 : _GEN_21; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_23 = 5'h17 == io_in_0_bits_ctrl_rfSrc1 ? rf_23 : _GEN_22; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_24 = 5'h18 == io_in_0_bits_ctrl_rfSrc1 ? rf_24 : _GEN_23; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_25 = 5'h19 == io_in_0_bits_ctrl_rfSrc1 ? rf_25 : _GEN_24; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_26 = 5'h1a == io_in_0_bits_ctrl_rfSrc1 ? rf_26 : _GEN_25; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_27 = 5'h1b == io_in_0_bits_ctrl_rfSrc1 ? rf_27 : _GEN_26; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_28 = 5'h1c == io_in_0_bits_ctrl_rfSrc1 ? rf_28 : _GEN_27; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_29 = 5'h1d == io_in_0_bits_ctrl_rfSrc1 ? rf_29 : _GEN_28; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_30 = 5'h1e == io_in_0_bits_ctrl_rfSrc1 ? rf_30 : _GEN_29; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_31 = 5'h1f == io_in_0_bits_ctrl_rfSrc1 ? rf_31 : _GEN_30; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _io_out_bits_data_src1_T_11 = io_in_0_bits_ctrl_rfSrc1 == 5'h0 ? 64'h0 : _GEN_31; // @[src/main/scala/nutcore/RF.scala 32:36]
  wire [63:0] _io_out_bits_data_src1_T_12 = io_in_0_bits_ctrl_src1Type ? _io_out_bits_data_src1_T_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_13 = src1ForwardNextCycle ? io_forward_wb_rfData : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_14 = _io_out_bits_data_src1_T_4 ? io_wb_rfData : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_15 = _io_out_bits_data_src1_T_9 ? _io_out_bits_data_src1_T_11 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_16 = _io_out_bits_data_src1_T_12 | _io_out_bits_data_src1_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src1_T_17 = _io_out_bits_data_src1_T_16 | _io_out_bits_data_src1_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_out_bits_data_src2_T_1 = ~src2ForwardNextCycle; // @[src/main/scala/nutcore/backend/seq/ISU.scala 72:21]
  wire  _io_out_bits_data_src2_T_2 = src2Forward & ~src2ForwardNextCycle; // @[src/main/scala/nutcore/backend/seq/ISU.scala 72:18]
  wire  _io_out_bits_data_src2_T_7 = ~io_in_0_bits_ctrl_src2Type & _io_out_bits_data_src2_T_1 & ~src2Forward; // @[src/main/scala/nutcore/backend/seq/ISU.scala 73:77]
  wire [63:0] _GEN_33 = 5'h1 == io_in_0_bits_ctrl_rfSrc2 ? rf_1 : rf_0; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_34 = 5'h2 == io_in_0_bits_ctrl_rfSrc2 ? rf_2 : _GEN_33; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_35 = 5'h3 == io_in_0_bits_ctrl_rfSrc2 ? rf_3 : _GEN_34; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_36 = 5'h4 == io_in_0_bits_ctrl_rfSrc2 ? rf_4 : _GEN_35; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_37 = 5'h5 == io_in_0_bits_ctrl_rfSrc2 ? rf_5 : _GEN_36; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_38 = 5'h6 == io_in_0_bits_ctrl_rfSrc2 ? rf_6 : _GEN_37; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_39 = 5'h7 == io_in_0_bits_ctrl_rfSrc2 ? rf_7 : _GEN_38; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_40 = 5'h8 == io_in_0_bits_ctrl_rfSrc2 ? rf_8 : _GEN_39; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_41 = 5'h9 == io_in_0_bits_ctrl_rfSrc2 ? rf_9 : _GEN_40; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_42 = 5'ha == io_in_0_bits_ctrl_rfSrc2 ? rf_10 : _GEN_41; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_43 = 5'hb == io_in_0_bits_ctrl_rfSrc2 ? rf_11 : _GEN_42; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_44 = 5'hc == io_in_0_bits_ctrl_rfSrc2 ? rf_12 : _GEN_43; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_45 = 5'hd == io_in_0_bits_ctrl_rfSrc2 ? rf_13 : _GEN_44; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_46 = 5'he == io_in_0_bits_ctrl_rfSrc2 ? rf_14 : _GEN_45; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_47 = 5'hf == io_in_0_bits_ctrl_rfSrc2 ? rf_15 : _GEN_46; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_48 = 5'h10 == io_in_0_bits_ctrl_rfSrc2 ? rf_16 : _GEN_47; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_49 = 5'h11 == io_in_0_bits_ctrl_rfSrc2 ? rf_17 : _GEN_48; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_50 = 5'h12 == io_in_0_bits_ctrl_rfSrc2 ? rf_18 : _GEN_49; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_51 = 5'h13 == io_in_0_bits_ctrl_rfSrc2 ? rf_19 : _GEN_50; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_52 = 5'h14 == io_in_0_bits_ctrl_rfSrc2 ? rf_20 : _GEN_51; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_53 = 5'h15 == io_in_0_bits_ctrl_rfSrc2 ? rf_21 : _GEN_52; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_54 = 5'h16 == io_in_0_bits_ctrl_rfSrc2 ? rf_22 : _GEN_53; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_55 = 5'h17 == io_in_0_bits_ctrl_rfSrc2 ? rf_23 : _GEN_54; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_56 = 5'h18 == io_in_0_bits_ctrl_rfSrc2 ? rf_24 : _GEN_55; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_57 = 5'h19 == io_in_0_bits_ctrl_rfSrc2 ? rf_25 : _GEN_56; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_58 = 5'h1a == io_in_0_bits_ctrl_rfSrc2 ? rf_26 : _GEN_57; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_59 = 5'h1b == io_in_0_bits_ctrl_rfSrc2 ? rf_27 : _GEN_58; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_60 = 5'h1c == io_in_0_bits_ctrl_rfSrc2 ? rf_28 : _GEN_59; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_61 = 5'h1d == io_in_0_bits_ctrl_rfSrc2 ? rf_29 : _GEN_60; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_62 = 5'h1e == io_in_0_bits_ctrl_rfSrc2 ? rf_30 : _GEN_61; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _GEN_63 = 5'h1f == io_in_0_bits_ctrl_rfSrc2 ? rf_31 : _GEN_62; // @[src/main/scala/nutcore/RF.scala 32:{36,36}]
  wire [63:0] _io_out_bits_data_src2_T_9 = io_in_0_bits_ctrl_rfSrc2 == 5'h0 ? 64'h0 : _GEN_63; // @[src/main/scala/nutcore/RF.scala 32:36]
  wire [63:0] _io_out_bits_data_src2_T_10 = io_in_0_bits_ctrl_src2Type ? io_in_0_bits_data_imm : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_11 = src2ForwardNextCycle ? io_forward_wb_rfData : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_12 = _io_out_bits_data_src2_T_2 ? io_wb_rfData : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_13 = _io_out_bits_data_src2_T_7 ? _io_out_bits_data_src2_T_9 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_14 = _io_out_bits_data_src2_T_10 | _io_out_bits_data_src2_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_out_bits_data_src2_T_15 = _io_out_bits_data_src2_T_14 | _io_out_bits_data_src2_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _wbClearMask_T_3 = io_wb_rfDest != 5'h0 & io_wb_rfDest == io_forward_wb_rfDest & forwardRfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 41:100]
  wire [62:0] _wbClearMask_T_6 = 63'h1 << io_wb_rfDest; // @[src/main/scala/nutcore/RF.scala 39:39]
  wire [31:0] wbClearMask = io_wb_rfWen & ~_wbClearMask_T_3 ? _wbClearMask_T_6[31:0] : 32'h0; // @[src/main/scala/nutcore/backend/seq/ISU.scala 85:24]
  wire  _isuFireSetMask_T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [62:0] _isuFireSetMask_T_1 = 63'h1 << io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/RF.scala 39:39]
  wire [31:0] isuFireSetMask = _isuFireSetMask_T ? _isuFireSetMask_T_1[31:0] : 32'h0; // @[src/main/scala/nutcore/backend/seq/ISU.scala 87:27]
  wire [31:0] _busy_T_5 = ~wbClearMask; // @[src/main/scala/nutcore/RF.scala 45:26]
  wire [31:0] _busy_T_6 = busy & _busy_T_5; // @[src/main/scala/nutcore/RF.scala 45:24]
  wire [31:0] _busy_T_7 = _busy_T_6 | isuFireSetMask; // @[src/main/scala/nutcore/RF.scala 45:38]
  wire [31:0] _busy_T_9 = {_busy_T_7[31:1],1'h0}; // @[src/main/scala/nutcore/RF.scala 45:16]
  wire  _T_3 = io_in_0_valid & ~io_out_valid; // @[src/main/scala/nutcore/backend/seq/ISU.scala 97:40]
  wire  _T_6 = io_out_valid & ~_isuFireSetMask_T; // @[src/main/scala/nutcore/backend/seq/ISU.scala 98:38]
  wire  _T_7 = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [31:0] busy_p; // @[src/main/scala/nutcore/RF.scala 37:21]
  wire [31:0] busy_t = busy ^ busy_p; // @[src/main/scala/nutcore/RF.scala 37:21]
  wire  toggle_504_clock;
  wire  toggle_504_reset;
  wire [31:0] toggle_504_valid;
  reg [31:0] toggle_504_valid_reg;
  reg [63:0] rf_0_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_0_t = rf_0 ^ rf_0_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_536_clock;
  wire  toggle_536_reset;
  wire [63:0] toggle_536_valid;
  reg [63:0] toggle_536_valid_reg;
  reg [63:0] rf_1_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_1_t = rf_1 ^ rf_1_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_600_clock;
  wire  toggle_600_reset;
  wire [63:0] toggle_600_valid;
  reg [63:0] toggle_600_valid_reg;
  reg [63:0] rf_2_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_2_t = rf_2 ^ rf_2_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_664_clock;
  wire  toggle_664_reset;
  wire [63:0] toggle_664_valid;
  reg [63:0] toggle_664_valid_reg;
  reg [63:0] rf_3_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_3_t = rf_3 ^ rf_3_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_728_clock;
  wire  toggle_728_reset;
  wire [63:0] toggle_728_valid;
  reg [63:0] toggle_728_valid_reg;
  reg [63:0] rf_4_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_4_t = rf_4 ^ rf_4_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_792_clock;
  wire  toggle_792_reset;
  wire [63:0] toggle_792_valid;
  reg [63:0] toggle_792_valid_reg;
  reg [63:0] rf_5_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_5_t = rf_5 ^ rf_5_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_856_clock;
  wire  toggle_856_reset;
  wire [63:0] toggle_856_valid;
  reg [63:0] toggle_856_valid_reg;
  reg [63:0] rf_6_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_6_t = rf_6 ^ rf_6_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_920_clock;
  wire  toggle_920_reset;
  wire [63:0] toggle_920_valid;
  reg [63:0] toggle_920_valid_reg;
  reg [63:0] rf_7_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_7_t = rf_7 ^ rf_7_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_984_clock;
  wire  toggle_984_reset;
  wire [63:0] toggle_984_valid;
  reg [63:0] toggle_984_valid_reg;
  reg [63:0] rf_8_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_8_t = rf_8 ^ rf_8_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_1048_clock;
  wire  toggle_1048_reset;
  wire [63:0] toggle_1048_valid;
  reg [63:0] toggle_1048_valid_reg;
  reg [63:0] rf_9_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_9_t = rf_9 ^ rf_9_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_1112_clock;
  wire  toggle_1112_reset;
  wire [63:0] toggle_1112_valid;
  reg [63:0] toggle_1112_valid_reg;
  reg [63:0] rf_10_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_10_t = rf_10 ^ rf_10_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_1176_clock;
  wire  toggle_1176_reset;
  wire [63:0] toggle_1176_valid;
  reg [63:0] toggle_1176_valid_reg;
  reg [63:0] rf_11_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_11_t = rf_11 ^ rf_11_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_1240_clock;
  wire  toggle_1240_reset;
  wire [63:0] toggle_1240_valid;
  reg [63:0] toggle_1240_valid_reg;
  reg [63:0] rf_12_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_12_t = rf_12 ^ rf_12_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_1304_clock;
  wire  toggle_1304_reset;
  wire [63:0] toggle_1304_valid;
  reg [63:0] toggle_1304_valid_reg;
  reg [63:0] rf_13_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_13_t = rf_13 ^ rf_13_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_1368_clock;
  wire  toggle_1368_reset;
  wire [63:0] toggle_1368_valid;
  reg [63:0] toggle_1368_valid_reg;
  reg [63:0] rf_14_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_14_t = rf_14 ^ rf_14_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_1432_clock;
  wire  toggle_1432_reset;
  wire [63:0] toggle_1432_valid;
  reg [63:0] toggle_1432_valid_reg;
  reg [63:0] rf_15_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_15_t = rf_15 ^ rf_15_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_1496_clock;
  wire  toggle_1496_reset;
  wire [63:0] toggle_1496_valid;
  reg [63:0] toggle_1496_valid_reg;
  reg [63:0] rf_16_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_16_t = rf_16 ^ rf_16_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_1560_clock;
  wire  toggle_1560_reset;
  wire [63:0] toggle_1560_valid;
  reg [63:0] toggle_1560_valid_reg;
  reg [63:0] rf_17_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_17_t = rf_17 ^ rf_17_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_1624_clock;
  wire  toggle_1624_reset;
  wire [63:0] toggle_1624_valid;
  reg [63:0] toggle_1624_valid_reg;
  reg [63:0] rf_18_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_18_t = rf_18 ^ rf_18_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_1688_clock;
  wire  toggle_1688_reset;
  wire [63:0] toggle_1688_valid;
  reg [63:0] toggle_1688_valid_reg;
  reg [63:0] rf_19_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_19_t = rf_19 ^ rf_19_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_1752_clock;
  wire  toggle_1752_reset;
  wire [63:0] toggle_1752_valid;
  reg [63:0] toggle_1752_valid_reg;
  reg [63:0] rf_20_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_20_t = rf_20 ^ rf_20_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_1816_clock;
  wire  toggle_1816_reset;
  wire [63:0] toggle_1816_valid;
  reg [63:0] toggle_1816_valid_reg;
  reg [63:0] rf_21_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_21_t = rf_21 ^ rf_21_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_1880_clock;
  wire  toggle_1880_reset;
  wire [63:0] toggle_1880_valid;
  reg [63:0] toggle_1880_valid_reg;
  reg [63:0] rf_22_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_22_t = rf_22 ^ rf_22_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_1944_clock;
  wire  toggle_1944_reset;
  wire [63:0] toggle_1944_valid;
  reg [63:0] toggle_1944_valid_reg;
  reg [63:0] rf_23_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_23_t = rf_23 ^ rf_23_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_2008_clock;
  wire  toggle_2008_reset;
  wire [63:0] toggle_2008_valid;
  reg [63:0] toggle_2008_valid_reg;
  reg [63:0] rf_24_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_24_t = rf_24 ^ rf_24_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_2072_clock;
  wire  toggle_2072_reset;
  wire [63:0] toggle_2072_valid;
  reg [63:0] toggle_2072_valid_reg;
  reg [63:0] rf_25_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_25_t = rf_25 ^ rf_25_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_2136_clock;
  wire  toggle_2136_reset;
  wire [63:0] toggle_2136_valid;
  reg [63:0] toggle_2136_valid_reg;
  reg [63:0] rf_26_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_26_t = rf_26 ^ rf_26_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_2200_clock;
  wire  toggle_2200_reset;
  wire [63:0] toggle_2200_valid;
  reg [63:0] toggle_2200_valid_reg;
  reg [63:0] rf_27_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_27_t = rf_27 ^ rf_27_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_2264_clock;
  wire  toggle_2264_reset;
  wire [63:0] toggle_2264_valid;
  reg [63:0] toggle_2264_valid_reg;
  reg [63:0] rf_28_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_28_t = rf_28 ^ rf_28_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_2328_clock;
  wire  toggle_2328_reset;
  wire [63:0] toggle_2328_valid;
  reg [63:0] toggle_2328_valid_reg;
  reg [63:0] rf_29_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_29_t = rf_29 ^ rf_29_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_2392_clock;
  wire  toggle_2392_reset;
  wire [63:0] toggle_2392_valid;
  reg [63:0] toggle_2392_valid_reg;
  reg [63:0] rf_30_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_30_t = rf_30 ^ rf_30_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_2456_clock;
  wire  toggle_2456_reset;
  wire [63:0] toggle_2456_valid;
  reg [63:0] toggle_2456_valid_reg;
  reg [63:0] rf_31_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire [63:0] rf_31_t = rf_31 ^ rf_31_p; // @[src/main/scala/nutcore/RF.scala 31:19]
  wire  toggle_2520_clock;
  wire  toggle_2520_reset;
  wire [63:0] toggle_2520_valid;
  reg [63:0] toggle_2520_valid_reg;
  DummyDPICWrapper difftest_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_clock),
    .reset(difftest_module_reset),
    .io_bits_value_1(difftest_module_io_bits_value_1),
    .io_bits_value_2(difftest_module_io_bits_value_2),
    .io_bits_value_3(difftest_module_io_bits_value_3),
    .io_bits_value_4(difftest_module_io_bits_value_4),
    .io_bits_value_5(difftest_module_io_bits_value_5),
    .io_bits_value_6(difftest_module_io_bits_value_6),
    .io_bits_value_7(difftest_module_io_bits_value_7),
    .io_bits_value_8(difftest_module_io_bits_value_8),
    .io_bits_value_9(difftest_module_io_bits_value_9),
    .io_bits_value_10(difftest_module_io_bits_value_10),
    .io_bits_value_11(difftest_module_io_bits_value_11),
    .io_bits_value_12(difftest_module_io_bits_value_12),
    .io_bits_value_13(difftest_module_io_bits_value_13),
    .io_bits_value_14(difftest_module_io_bits_value_14),
    .io_bits_value_15(difftest_module_io_bits_value_15),
    .io_bits_value_16(difftest_module_io_bits_value_16),
    .io_bits_value_17(difftest_module_io_bits_value_17),
    .io_bits_value_18(difftest_module_io_bits_value_18),
    .io_bits_value_19(difftest_module_io_bits_value_19),
    .io_bits_value_20(difftest_module_io_bits_value_20),
    .io_bits_value_21(difftest_module_io_bits_value_21),
    .io_bits_value_22(difftest_module_io_bits_value_22),
    .io_bits_value_23(difftest_module_io_bits_value_23),
    .io_bits_value_24(difftest_module_io_bits_value_24),
    .io_bits_value_25(difftest_module_io_bits_value_25),
    .io_bits_value_26(difftest_module_io_bits_value_26),
    .io_bits_value_27(difftest_module_io_bits_value_27),
    .io_bits_value_28(difftest_module_io_bits_value_28),
    .io_bits_value_29(difftest_module_io_bits_value_29),
    .io_bits_value_30(difftest_module_io_bits_value_30),
    .io_bits_value_31(difftest_module_io_bits_value_31)
  );
  GEN_w32_toggle #(.COVER_INDEX(504)) toggle_504 (
    .clock(toggle_504_clock),
    .reset(toggle_504_reset),
    .valid(toggle_504_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(536)) toggle_536 (
    .clock(toggle_536_clock),
    .reset(toggle_536_reset),
    .valid(toggle_536_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(600)) toggle_600 (
    .clock(toggle_600_clock),
    .reset(toggle_600_reset),
    .valid(toggle_600_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(664)) toggle_664 (
    .clock(toggle_664_clock),
    .reset(toggle_664_reset),
    .valid(toggle_664_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(728)) toggle_728 (
    .clock(toggle_728_clock),
    .reset(toggle_728_reset),
    .valid(toggle_728_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(792)) toggle_792 (
    .clock(toggle_792_clock),
    .reset(toggle_792_reset),
    .valid(toggle_792_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(856)) toggle_856 (
    .clock(toggle_856_clock),
    .reset(toggle_856_reset),
    .valid(toggle_856_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(920)) toggle_920 (
    .clock(toggle_920_clock),
    .reset(toggle_920_reset),
    .valid(toggle_920_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(984)) toggle_984 (
    .clock(toggle_984_clock),
    .reset(toggle_984_reset),
    .valid(toggle_984_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(1048)) toggle_1048 (
    .clock(toggle_1048_clock),
    .reset(toggle_1048_reset),
    .valid(toggle_1048_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(1112)) toggle_1112 (
    .clock(toggle_1112_clock),
    .reset(toggle_1112_reset),
    .valid(toggle_1112_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(1176)) toggle_1176 (
    .clock(toggle_1176_clock),
    .reset(toggle_1176_reset),
    .valid(toggle_1176_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(1240)) toggle_1240 (
    .clock(toggle_1240_clock),
    .reset(toggle_1240_reset),
    .valid(toggle_1240_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(1304)) toggle_1304 (
    .clock(toggle_1304_clock),
    .reset(toggle_1304_reset),
    .valid(toggle_1304_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(1368)) toggle_1368 (
    .clock(toggle_1368_clock),
    .reset(toggle_1368_reset),
    .valid(toggle_1368_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(1432)) toggle_1432 (
    .clock(toggle_1432_clock),
    .reset(toggle_1432_reset),
    .valid(toggle_1432_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(1496)) toggle_1496 (
    .clock(toggle_1496_clock),
    .reset(toggle_1496_reset),
    .valid(toggle_1496_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(1560)) toggle_1560 (
    .clock(toggle_1560_clock),
    .reset(toggle_1560_reset),
    .valid(toggle_1560_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(1624)) toggle_1624 (
    .clock(toggle_1624_clock),
    .reset(toggle_1624_reset),
    .valid(toggle_1624_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(1688)) toggle_1688 (
    .clock(toggle_1688_clock),
    .reset(toggle_1688_reset),
    .valid(toggle_1688_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(1752)) toggle_1752 (
    .clock(toggle_1752_clock),
    .reset(toggle_1752_reset),
    .valid(toggle_1752_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(1816)) toggle_1816 (
    .clock(toggle_1816_clock),
    .reset(toggle_1816_reset),
    .valid(toggle_1816_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(1880)) toggle_1880 (
    .clock(toggle_1880_clock),
    .reset(toggle_1880_reset),
    .valid(toggle_1880_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(1944)) toggle_1944 (
    .clock(toggle_1944_clock),
    .reset(toggle_1944_reset),
    .valid(toggle_1944_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(2008)) toggle_2008 (
    .clock(toggle_2008_clock),
    .reset(toggle_2008_reset),
    .valid(toggle_2008_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(2072)) toggle_2072 (
    .clock(toggle_2072_clock),
    .reset(toggle_2072_reset),
    .valid(toggle_2072_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(2136)) toggle_2136 (
    .clock(toggle_2136_clock),
    .reset(toggle_2136_reset),
    .valid(toggle_2136_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(2200)) toggle_2200 (
    .clock(toggle_2200_clock),
    .reset(toggle_2200_reset),
    .valid(toggle_2200_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(2264)) toggle_2264 (
    .clock(toggle_2264_clock),
    .reset(toggle_2264_reset),
    .valid(toggle_2264_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(2328)) toggle_2328 (
    .clock(toggle_2328_clock),
    .reset(toggle_2328_reset),
    .valid(toggle_2328_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(2392)) toggle_2392 (
    .clock(toggle_2392_clock),
    .reset(toggle_2392_reset),
    .valid(toggle_2392_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(2456)) toggle_2456 (
    .clock(toggle_2456_clock),
    .reset(toggle_2456_reset),
    .valid(toggle_2456_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(2520)) toggle_2520 (
    .clock(toggle_2520_clock),
    .reset(toggle_2520_reset),
    .valid(toggle_2520_valid)
  );
  assign io_in_0_ready = ~io_in_0_valid | _isuFireSetMask_T; // @[src/main/scala/nutcore/backend/seq/ISU.scala 91:37]
  assign io_out_valid = io_in_0_valid & src1Ready & src2Ready; // @[src/main/scala/nutcore/backend/seq/ISU.scala 58:47]
  assign io_out_bits_cf_instr = io_in_0_bits_cf_instr; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_pc = io_in_0_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_pnpc = io_in_0_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_exceptionVec_1 = io_in_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_exceptionVec_2 = io_in_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_exceptionVec_12 = io_in_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_1 = io_in_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_3 = io_in_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_5 = io_in_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_7 = io_in_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_9 = io_in_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_intrVec_11 = io_in_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_brIdx = io_in_0_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_cf_crossBoundaryFault = io_in_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/backend/seq/ISU.scala 77:18]
  assign io_out_bits_ctrl_fuType = io_in_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_fuOpType = io_in_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_rfWen = io_in_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_rfDest = io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_ctrl_isNutCoreTrap = io_in_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/seq/ISU.scala 78:20]
  assign io_out_bits_data_src1 = _io_out_bits_data_src1_T_17 | _io_out_bits_data_src1_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_bits_data_src2 = _io_out_bits_data_src2_T_15 | _io_out_bits_data_src2_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_bits_data_imm = io_in_0_bits_data_imm; // @[src/main/scala/nutcore/backend/seq/ISU.scala 75:25]
  assign difftest_module_clock = clock;
  assign difftest_module_reset = reset;
  assign difftest_module_io_bits_value_1 = rf_1; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_2 = rf_2; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_3 = rf_3; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_4 = rf_4; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_5 = rf_5; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_6 = rf_6; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_7 = rf_7; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_8 = rf_8; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_9 = rf_9; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_10 = rf_10; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_11 = rf_11; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_12 = rf_12; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_13 = rf_13; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_14 = rf_14; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_15 = rf_15; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_16 = rf_16; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_17 = rf_17; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_18 = rf_18; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_19 = rf_19; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_20 = rf_20; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_21 = rf_21; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_22 = rf_22; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_23 = rf_23; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_24 = rf_24; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_25 = rf_25; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_26 = rf_26; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_27 = rf_27; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_28 = rf_28; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_29 = rf_29; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_30 = rf_30; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign difftest_module_io_bits_value_31 = rf_31; // @[src/main/scala/nutcore/RF.scala 32:36]
  assign toggle_504_clock = clock;
  assign toggle_504_reset = reset;
  assign toggle_504_valid = busy ^ toggle_504_valid_reg;
  assign toggle_536_clock = clock;
  assign toggle_536_reset = reset;
  assign toggle_536_valid = rf_0 ^ toggle_536_valid_reg;
  assign toggle_600_clock = clock;
  assign toggle_600_reset = reset;
  assign toggle_600_valid = rf_1 ^ toggle_600_valid_reg;
  assign toggle_664_clock = clock;
  assign toggle_664_reset = reset;
  assign toggle_664_valid = rf_2 ^ toggle_664_valid_reg;
  assign toggle_728_clock = clock;
  assign toggle_728_reset = reset;
  assign toggle_728_valid = rf_3 ^ toggle_728_valid_reg;
  assign toggle_792_clock = clock;
  assign toggle_792_reset = reset;
  assign toggle_792_valid = rf_4 ^ toggle_792_valid_reg;
  assign toggle_856_clock = clock;
  assign toggle_856_reset = reset;
  assign toggle_856_valid = rf_5 ^ toggle_856_valid_reg;
  assign toggle_920_clock = clock;
  assign toggle_920_reset = reset;
  assign toggle_920_valid = rf_6 ^ toggle_920_valid_reg;
  assign toggle_984_clock = clock;
  assign toggle_984_reset = reset;
  assign toggle_984_valid = rf_7 ^ toggle_984_valid_reg;
  assign toggle_1048_clock = clock;
  assign toggle_1048_reset = reset;
  assign toggle_1048_valid = rf_8 ^ toggle_1048_valid_reg;
  assign toggle_1112_clock = clock;
  assign toggle_1112_reset = reset;
  assign toggle_1112_valid = rf_9 ^ toggle_1112_valid_reg;
  assign toggle_1176_clock = clock;
  assign toggle_1176_reset = reset;
  assign toggle_1176_valid = rf_10 ^ toggle_1176_valid_reg;
  assign toggle_1240_clock = clock;
  assign toggle_1240_reset = reset;
  assign toggle_1240_valid = rf_11 ^ toggle_1240_valid_reg;
  assign toggle_1304_clock = clock;
  assign toggle_1304_reset = reset;
  assign toggle_1304_valid = rf_12 ^ toggle_1304_valid_reg;
  assign toggle_1368_clock = clock;
  assign toggle_1368_reset = reset;
  assign toggle_1368_valid = rf_13 ^ toggle_1368_valid_reg;
  assign toggle_1432_clock = clock;
  assign toggle_1432_reset = reset;
  assign toggle_1432_valid = rf_14 ^ toggle_1432_valid_reg;
  assign toggle_1496_clock = clock;
  assign toggle_1496_reset = reset;
  assign toggle_1496_valid = rf_15 ^ toggle_1496_valid_reg;
  assign toggle_1560_clock = clock;
  assign toggle_1560_reset = reset;
  assign toggle_1560_valid = rf_16 ^ toggle_1560_valid_reg;
  assign toggle_1624_clock = clock;
  assign toggle_1624_reset = reset;
  assign toggle_1624_valid = rf_17 ^ toggle_1624_valid_reg;
  assign toggle_1688_clock = clock;
  assign toggle_1688_reset = reset;
  assign toggle_1688_valid = rf_18 ^ toggle_1688_valid_reg;
  assign toggle_1752_clock = clock;
  assign toggle_1752_reset = reset;
  assign toggle_1752_valid = rf_19 ^ toggle_1752_valid_reg;
  assign toggle_1816_clock = clock;
  assign toggle_1816_reset = reset;
  assign toggle_1816_valid = rf_20 ^ toggle_1816_valid_reg;
  assign toggle_1880_clock = clock;
  assign toggle_1880_reset = reset;
  assign toggle_1880_valid = rf_21 ^ toggle_1880_valid_reg;
  assign toggle_1944_clock = clock;
  assign toggle_1944_reset = reset;
  assign toggle_1944_valid = rf_22 ^ toggle_1944_valid_reg;
  assign toggle_2008_clock = clock;
  assign toggle_2008_reset = reset;
  assign toggle_2008_valid = rf_23 ^ toggle_2008_valid_reg;
  assign toggle_2072_clock = clock;
  assign toggle_2072_reset = reset;
  assign toggle_2072_valid = rf_24 ^ toggle_2072_valid_reg;
  assign toggle_2136_clock = clock;
  assign toggle_2136_reset = reset;
  assign toggle_2136_valid = rf_25 ^ toggle_2136_valid_reg;
  assign toggle_2200_clock = clock;
  assign toggle_2200_reset = reset;
  assign toggle_2200_valid = rf_26 ^ toggle_2200_valid_reg;
  assign toggle_2264_clock = clock;
  assign toggle_2264_reset = reset;
  assign toggle_2264_valid = rf_27 ^ toggle_2264_valid_reg;
  assign toggle_2328_clock = clock;
  assign toggle_2328_reset = reset;
  assign toggle_2328_valid = rf_28 ^ toggle_2328_valid_reg;
  assign toggle_2392_clock = clock;
  assign toggle_2392_reset = reset;
  assign toggle_2392_valid = rf_29 ^ toggle_2392_valid_reg;
  assign toggle_2456_clock = clock;
  assign toggle_2456_reset = reset;
  assign toggle_2456_valid = rf_30 ^ toggle_2456_valid_reg;
  assign toggle_2520_clock = clock;
  assign toggle_2520_reset = reset;
  assign toggle_2520_valid = rf_31 ^ toggle_2520_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 37:21]
      busy <= 32'h0; // @[src/main/scala/nutcore/RF.scala 37:21]
    end else if (io_flush) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 88:19]
      busy <= 32'h0; // @[src/main/scala/nutcore/RF.scala 45:10]
    end else begin
      busy <= _busy_T_9; // @[src/main/scala/nutcore/RF.scala 45:10]
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_0 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h0 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_0 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_1 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_1 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_2 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h2 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_2 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_3 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h3 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_3 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_4 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h4 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_4 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_5 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h5 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_5 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_6 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h6 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_6 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_7 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h7 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_7 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_8 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h8 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_8 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_9 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h9 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_9 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_10 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'ha == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_10 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_11 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'hb == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_11 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_12 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'hc == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_12 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_13 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'hd == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_13 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_14 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'he == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_14 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_15 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'hf == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_15 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_16 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h10 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_16 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_17 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h11 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_17 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_18 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h12 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_18 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_19 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h13 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_19 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_20 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h14 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_20 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_21 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h15 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_21 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_22 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h16 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_22 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_23 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h17 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_23 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_24 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h18 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_24 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_25 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h19 == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_25 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_26 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1a == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_26 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_27 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1b == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_27 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_28 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1c == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_28 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_29 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1d == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_29 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_30 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1e == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_30 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/RF.scala 31:19]
      rf_31 <= 64'h0; // @[src/main/scala/nutcore/RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[src/main/scala/nutcore/backend/seq/ISU.scala 83:22]
      if (5'h1f == io_wb_rfDest) begin // @[src/main/scala/nutcore/RF.scala 33:50]
        rf_31 <= io_wb_rfData; // @[src/main/scala/nutcore/RF.scala 33:50]
      end
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    busy_p <= busy; // @[src/main/scala/nutcore/RF.scala 37:21]
    toggle_504_valid_reg <= busy;
    rf_0_p <= rf_0; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_536_valid_reg <= rf_0;
    rf_1_p <= rf_1; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_600_valid_reg <= rf_1;
    rf_2_p <= rf_2; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_664_valid_reg <= rf_2;
    rf_3_p <= rf_3; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_728_valid_reg <= rf_3;
    rf_4_p <= rf_4; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_792_valid_reg <= rf_4;
    rf_5_p <= rf_5; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_856_valid_reg <= rf_5;
    rf_6_p <= rf_6; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_920_valid_reg <= rf_6;
    rf_7_p <= rf_7; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_984_valid_reg <= rf_7;
    rf_8_p <= rf_8; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_1048_valid_reg <= rf_8;
    rf_9_p <= rf_9; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_1112_valid_reg <= rf_9;
    rf_10_p <= rf_10; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_1176_valid_reg <= rf_10;
    rf_11_p <= rf_11; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_1240_valid_reg <= rf_11;
    rf_12_p <= rf_12; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_1304_valid_reg <= rf_12;
    rf_13_p <= rf_13; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_1368_valid_reg <= rf_13;
    rf_14_p <= rf_14; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_1432_valid_reg <= rf_14;
    rf_15_p <= rf_15; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_1496_valid_reg <= rf_15;
    rf_16_p <= rf_16; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_1560_valid_reg <= rf_16;
    rf_17_p <= rf_17; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_1624_valid_reg <= rf_17;
    rf_18_p <= rf_18; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_1688_valid_reg <= rf_18;
    rf_19_p <= rf_19; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_1752_valid_reg <= rf_19;
    rf_20_p <= rf_20; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_1816_valid_reg <= rf_20;
    rf_21_p <= rf_21; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_1880_valid_reg <= rf_21;
    rf_22_p <= rf_22; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_1944_valid_reg <= rf_22;
    rf_23_p <= rf_23; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_2008_valid_reg <= rf_23;
    rf_24_p <= rf_24; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_2072_valid_reg <= rf_24;
    rf_25_p <= rf_25; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_2136_valid_reg <= rf_25;
    rf_26_p <= rf_26; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_2200_valid_reg <= rf_26;
    rf_27_p <= rf_27; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_2264_valid_reg <= rf_27;
    rf_28_p <= rf_28; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_2328_valid_reg <= rf_28;
    rf_29_p <= rf_29; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_2392_valid_reg <= rf_29;
    rf_30_p <= rf_30; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_2456_valid_reg <= rf_30;
    rf_31_p <= rf_31; // @[src/main/scala/nutcore/RF.scala 31:19]
    toggle_2520_valid_reg <= rf_31;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  busy = _RAND_0[31:0];
  _RAND_1 = {2{`RANDOM}};
  rf_0 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  rf_1 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  rf_2 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  rf_3 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  rf_4 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  rf_5 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  rf_6 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  rf_7 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  rf_8 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  rf_9 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  rf_10 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  rf_11 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  rf_12 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  rf_13 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  rf_14 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  rf_15 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  rf_16 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  rf_17 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  rf_18 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  rf_19 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  rf_20 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  rf_21 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  rf_22 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  rf_23 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  rf_24 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  rf_25 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  rf_26 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  rf_27 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  rf_28 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  rf_29 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  rf_30 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  rf_31 = _RAND_32[63:0];
  _RAND_33 = {1{`RANDOM}};
  busy_p = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  toggle_504_valid_reg = _RAND_34[31:0];
  _RAND_35 = {2{`RANDOM}};
  rf_0_p = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  toggle_536_valid_reg = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  rf_1_p = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  toggle_600_valid_reg = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  rf_2_p = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  toggle_664_valid_reg = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  rf_3_p = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  toggle_728_valid_reg = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  rf_4_p = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  toggle_792_valid_reg = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  rf_5_p = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  toggle_856_valid_reg = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  rf_6_p = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  toggle_920_valid_reg = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  rf_7_p = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  toggle_984_valid_reg = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  rf_8_p = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  toggle_1048_valid_reg = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  rf_9_p = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  toggle_1112_valid_reg = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  rf_10_p = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  toggle_1176_valid_reg = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  rf_11_p = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  toggle_1240_valid_reg = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  rf_12_p = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  toggle_1304_valid_reg = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  rf_13_p = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  toggle_1368_valid_reg = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  rf_14_p = _RAND_63[63:0];
  _RAND_64 = {2{`RANDOM}};
  toggle_1432_valid_reg = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  rf_15_p = _RAND_65[63:0];
  _RAND_66 = {2{`RANDOM}};
  toggle_1496_valid_reg = _RAND_66[63:0];
  _RAND_67 = {2{`RANDOM}};
  rf_16_p = _RAND_67[63:0];
  _RAND_68 = {2{`RANDOM}};
  toggle_1560_valid_reg = _RAND_68[63:0];
  _RAND_69 = {2{`RANDOM}};
  rf_17_p = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  toggle_1624_valid_reg = _RAND_70[63:0];
  _RAND_71 = {2{`RANDOM}};
  rf_18_p = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  toggle_1688_valid_reg = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  rf_19_p = _RAND_73[63:0];
  _RAND_74 = {2{`RANDOM}};
  toggle_1752_valid_reg = _RAND_74[63:0];
  _RAND_75 = {2{`RANDOM}};
  rf_20_p = _RAND_75[63:0];
  _RAND_76 = {2{`RANDOM}};
  toggle_1816_valid_reg = _RAND_76[63:0];
  _RAND_77 = {2{`RANDOM}};
  rf_21_p = _RAND_77[63:0];
  _RAND_78 = {2{`RANDOM}};
  toggle_1880_valid_reg = _RAND_78[63:0];
  _RAND_79 = {2{`RANDOM}};
  rf_22_p = _RAND_79[63:0];
  _RAND_80 = {2{`RANDOM}};
  toggle_1944_valid_reg = _RAND_80[63:0];
  _RAND_81 = {2{`RANDOM}};
  rf_23_p = _RAND_81[63:0];
  _RAND_82 = {2{`RANDOM}};
  toggle_2008_valid_reg = _RAND_82[63:0];
  _RAND_83 = {2{`RANDOM}};
  rf_24_p = _RAND_83[63:0];
  _RAND_84 = {2{`RANDOM}};
  toggle_2072_valid_reg = _RAND_84[63:0];
  _RAND_85 = {2{`RANDOM}};
  rf_25_p = _RAND_85[63:0];
  _RAND_86 = {2{`RANDOM}};
  toggle_2136_valid_reg = _RAND_86[63:0];
  _RAND_87 = {2{`RANDOM}};
  rf_26_p = _RAND_87[63:0];
  _RAND_88 = {2{`RANDOM}};
  toggle_2200_valid_reg = _RAND_88[63:0];
  _RAND_89 = {2{`RANDOM}};
  rf_27_p = _RAND_89[63:0];
  _RAND_90 = {2{`RANDOM}};
  toggle_2264_valid_reg = _RAND_90[63:0];
  _RAND_91 = {2{`RANDOM}};
  rf_28_p = _RAND_91[63:0];
  _RAND_92 = {2{`RANDOM}};
  toggle_2328_valid_reg = _RAND_92[63:0];
  _RAND_93 = {2{`RANDOM}};
  rf_29_p = _RAND_93[63:0];
  _RAND_94 = {2{`RANDOM}};
  toggle_2392_valid_reg = _RAND_94[63:0];
  _RAND_95 = {2{`RANDOM}};
  rf_30_p = _RAND_95[63:0];
  _RAND_96 = {2{`RANDOM}};
  toggle_2456_valid_reg = _RAND_96[63:0];
  _RAND_97 = {2{`RANDOM}};
  rf_31_p = _RAND_97[63:0];
  _RAND_98 = {2{`RANDOM}};
  toggle_2520_valid_reg = _RAND_98[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(busy_t[0]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[1]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[2]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[3]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[4]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[5]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[6]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[7]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[8]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[9]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[10]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[11]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[12]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[13]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[14]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[15]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[16]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[17]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[18]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[19]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[20]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[21]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[22]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[23]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[24]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[25]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[26]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[27]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[28]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[29]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[30]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(busy_t[31]); // @[src/main/scala/nutcore/RF.scala 37:21]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_0_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_1_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_2_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_3_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_4_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_5_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_6_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_7_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_8_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_9_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_10_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_11_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_12_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_13_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_14_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_15_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_16_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_17_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_18_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_19_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_20_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_21_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_22_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_23_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_24_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_25_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_26_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_27_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_28_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_29_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_30_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[0]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[1]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[2]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[3]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[4]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[5]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[6]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[7]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[8]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[9]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[10]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[11]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[12]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[13]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[14]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[15]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[16]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[17]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[18]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[19]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[20]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[21]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[22]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[23]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[24]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[25]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[26]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[27]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[28]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[29]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[30]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[31]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[32]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[33]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[34]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[35]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[36]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[37]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[38]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[39]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[40]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[41]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[42]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[43]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[44]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[45]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[46]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[47]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[48]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[49]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[50]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[51]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[52]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[53]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[54]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[55]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[56]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[57]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[58]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[59]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[60]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[61]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[62]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
    //
    if (enToggle_past) begin
      cover(rf_31_t[63]); // @[src/main/scala/nutcore/RF.scala 31:19]
    end
  end
endmodule
module ALU(
  input         clock,
  input         reset,
  input         io_in_valid, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [63:0] io_in_bits_src1, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [63:0] io_in_bits_src2, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [6:0]  io_in_bits_func, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output [63:0] io_out_bits, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [63:0] io_cfIn_instr, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [38:0] io_cfIn_pc, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [38:0] io_cfIn_pnpc, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [3:0]  io_cfIn_brIdx, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output [38:0] io_redirect_target, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output        io_redirect_valid, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input  [63:0] io_offset, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input         io_iVmEnable, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  input         io_jumpIsIllegal_ready, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output        io_jumpIsIllegal_valid, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output [63:0] io_jumpIsIllegal_bits, // @[src/main/scala/nutcore/backend/fu/ALU.scala 78:14]
  output        REG_0_valid,
  output [38:0] REG_0_pc,
  output        REG_0_isMissPredict,
  output [38:0] REG_0_actualTarget,
  output [6:0]  REG_0_fuOpType,
  output [1:0]  REG_0_btbType,
  output        REG_0_isRVC
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
`endif // RANDOMIZE_REG_INIT
  wire  isAdderSub = ~io_in_bits_func[6]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 89:20]
  wire [63:0] _adderRes_T = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[src/main/scala/nutcore/backend/fu/ALU.scala 90:39]
  wire [63:0] _adderRes_T_1 = io_in_bits_src2 ^ _adderRes_T; // @[src/main/scala/nutcore/backend/fu/ALU.scala 90:33]
  wire [64:0] _adderRes_T_2 = io_in_bits_src1 + _adderRes_T_1; // @[src/main/scala/nutcore/backend/fu/ALU.scala 90:24]
  wire [64:0] _GEN_12 = {{64'd0}, isAdderSub}; // @[src/main/scala/nutcore/backend/fu/ALU.scala 90:60]
  wire [64:0] adderRes = _adderRes_T_2 + _GEN_12; // @[src/main/scala/nutcore/backend/fu/ALU.scala 90:60]
  wire [63:0] xorRes = io_in_bits_src1 ^ io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 91:21]
  wire  sltu = ~adderRes[64]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 92:14]
  wire  slt = xorRes[63] ^ sltu; // @[src/main/scala/nutcore/backend/fu/ALU.scala 93:28]
  wire [63:0] _shsrc1_T_2 = {32'h0,io_in_bits_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  shsrc1_signBit = io_in_bits_src1[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _shsrc1_T_4 = shsrc1_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _shsrc1_T_5 = {_shsrc1_T_4,io_in_bits_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _shsrc1_T_7 = 7'h25 == io_in_bits_func ? _shsrc1_T_2 : io_in_bits_src1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [63:0] shsrc1 = 7'h2d == io_in_bits_func ? _shsrc1_T_5 : _shsrc1_T_7; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [5:0] shamt = io_in_bits_func[5] ? {{1'd0}, io_in_bits_src2[4:0]} : io_in_bits_src2[5:0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 99:18]
  wire [126:0] _GEN_15 = {{63'd0}, shsrc1}; // @[src/main/scala/nutcore/backend/fu/ALU.scala 101:33]
  wire [126:0] _res_T_1 = _GEN_15 << shamt; // @[src/main/scala/nutcore/backend/fu/ALU.scala 101:33]
  wire [63:0] _res_T_3 = {63'h0,slt}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _res_T_4 = {63'h0,sltu}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _res_T_5 = shsrc1 >> shamt; // @[src/main/scala/nutcore/backend/fu/ALU.scala 105:32]
  wire [63:0] _res_T_6 = io_in_bits_src1 | io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 106:30]
  wire [63:0] _res_T_7 = io_in_bits_src1 & io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 107:30]
  wire [63:0] _res_T_8 = 7'h2d == io_in_bits_func ? _shsrc1_T_5 : _shsrc1_T_7; // @[src/main/scala/nutcore/backend/fu/ALU.scala 108:32]
  wire [63:0] _res_T_10 = $signed(_res_T_8) >>> shamt; // @[src/main/scala/nutcore/backend/fu/ALU.scala 108:49]
  wire [64:0] _res_T_12 = 4'h1 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_1[63:0]} : adderRes; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_14 = 4'h2 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_3} : _res_T_12; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_16 = 4'h3 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_4} : _res_T_14; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_18 = 4'h4 == io_in_bits_func[3:0] ? {{1'd0}, xorRes} : _res_T_16; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_20 = 4'h5 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_5} : _res_T_18; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_22 = 4'h6 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_6} : _res_T_20; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_24 = 4'h7 == io_in_bits_func[3:0] ? {{1'd0}, _res_T_7} : _res_T_22; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] res = 4'hd == io_in_bits_func[3:0] ? {{1'd0}, _res_T_10} : _res_T_24; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  aluRes_signBit = res[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _aluRes_T_2 = aluRes_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _aluRes_T_3 = {_aluRes_T_2,res[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [64:0] aluRes = io_in_bits_func[5] ? {{1'd0}, _aluRes_T_3} : res; // @[src/main/scala/nutcore/backend/fu/ALU.scala 110:19]
  wire  _T_1 = ~(|xorRes); // @[src/main/scala/nutcore/backend/fu/ALU.scala 113:48]
  wire  isBranch = ~io_in_bits_func[3]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 63:30]
  wire  isBru = io_in_bits_func[4]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 62:31]
  wire  _taken_T_1 = 2'h0 == io_in_bits_func[2:1]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _taken_T_2 = 2'h2 == io_in_bits_func[2:1]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _taken_T_3 = 2'h3 == io_in_bits_func[2:1]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _taken_T_8 = _taken_T_1 & _T_1 | _taken_T_2 & slt | _taken_T_3 & sltu; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  taken = _taken_T_8 ^ io_in_bits_func[0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 120:72]
  wire  target_signBit = io_cfIn_pc[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _target_T = target_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _target_T_1 = {_target_T,io_cfIn_pc}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _target_T_3 = _target_T_1 + io_offset; // @[src/main/scala/nutcore/backend/fu/ALU.scala 121:56]
  wire [63:0] _target_T_5 = {adderRes[63:1],1'h0}; // @[src/main/scala/nutcore/backend/fu/ALU.scala 121:72]
  wire [63:0] target = isBranch ? _target_T_3 : _target_T_5; // @[src/main/scala/nutcore/backend/fu/ALU.scala 121:19]
  wire  _predictWrong_T_1 = ~taken & isBranch; // @[src/main/scala/nutcore/backend/fu/ALU.scala 122:33]
  wire  predictWrong = ~taken & isBranch ? io_cfIn_brIdx[0] : ~io_cfIn_brIdx[0] | io_redirect_target != io_cfIn_pnpc; // @[src/main/scala/nutcore/backend/fu/ALU.scala 122:25]
  wire  isRVC = io_cfIn_instr[1:0] != 2'h3; // @[src/main/scala/nutcore/backend/fu/ALU.scala 123:35]
  wire  _T_12 = ~isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 125:55]
  wire [38:0] _io_redirect_target_T_3 = io_cfIn_pc + 39'h2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 126:71]
  wire [38:0] _io_redirect_target_T_5 = io_cfIn_pc + 39'h4; // @[src/main/scala/nutcore/backend/fu/ALU.scala 126:89]
  wire [38:0] _io_redirect_target_T_6 = isRVC ? _io_redirect_target_T_3 : _io_redirect_target_T_5; // @[src/main/scala/nutcore/backend/fu/ALU.scala 126:52]
  wire [63:0] _io_redirect_target_T_7 = _predictWrong_T_1 ? {{25'd0}, _io_redirect_target_T_6} : target; // @[src/main/scala/nutcore/backend/fu/ALU.scala 126:28]
  wire  _io_redirect_valid_T = io_in_valid & isBru; // @[src/main/scala/nutcore/backend/fu/ALU.scala 128:30]
  wire  _io_redirect_valid_T_1 = io_in_valid & isBru & predictWrong; // @[src/main/scala/nutcore/backend/fu/ALU.scala 128:39]
  wire [63:0] _io_out_bits_T_4 = _target_T_1 + 64'h4; // @[src/main/scala/nutcore/backend/fu/ALU.scala 134:71]
  wire [63:0] _io_out_bits_T_8 = _target_T_1 + 64'h2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 134:108]
  wire [63:0] _io_out_bits_T_9 = _T_12 ? _io_out_bits_T_4 : _io_out_bits_T_8; // @[src/main/scala/nutcore/backend/fu/ALU.scala 134:32]
  wire [64:0] _io_out_bits_T_10 = isBru ? {{1'd0}, _io_out_bits_T_9} : aluRes; // @[src/main/scala/nutcore/backend/fu/ALU.scala 134:21]
  reg  hasIllegalJumpAddr; // @[src/main/scala/nutcore/backend/fu/ALU.scala 138:35]
  wire  addrNotLegal_signBit = target[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _addrNotLegal_T_1 = addrNotLegal_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _addrNotLegal_T_2 = {_addrNotLegal_T_1,target[38:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  addrNotLegal = io_iVmEnable ? target != _addrNotLegal_T_2 : |target[63:39]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 139:25]
  wire  isIllegalJumpAddr = io_redirect_valid & ~isBranch & addrNotLegal; // @[src/main/scala/nutcore/backend/fu/ALU.scala 140:58]
  wire  _T_15 = io_jumpIsIllegal_ready & io_jumpIsIllegal_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _GEN_0 = _T_15 ? 1'h0 : hasIllegalJumpAddr; // @[src/main/scala/nutcore/backend/fu/ALU.scala 143:38 144:24 138:35]
  wire  _GEN_1 = isIllegalJumpAddr | _GEN_0; // @[src/main/scala/nutcore/backend/fu/ALU.scala 141:28 142:24]
  reg [63:0] io_jumpIsIllegal_bits_r; // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
  wire  _T_21 = io_in_bits_func == 7'h58 | io_in_bits_func == 7'h5c; // @[src/main/scala/nutcore/backend/fu/ALU.scala 151:180]
  wire  _T_22 = io_in_bits_func == 7'h5a; // @[src/main/scala/nutcore/backend/fu/ALU.scala 151:214]
  wire  _T_23 = io_in_bits_func == 7'h5e; // @[src/main/scala/nutcore/backend/fu/ALU.scala 151:239]
  wire  _T_32 = 7'h5c == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _T_33 = 7'h5e == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _T_34 = 7'h58 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _T_35 = 7'h5a == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [1:0] _T_43 = _T_33 ? 2'h3 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _T_45 = _T_35 ? 2'h2 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _GEN_13 = {{1'd0}, _T_32}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _T_52 = _GEN_13 | _T_43; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _GEN_14 = {{1'd0}, _T_34}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _T_53 = _T_52 | _GEN_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  reg  REG_valid; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg [38:0] REG_pc; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg  REG_isMissPredict; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg [38:0] REG_actualTarget; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg  REG_actualTaken; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg [6:0] REG_fuOpType; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg [1:0] REG_btbType; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  reg  REG_isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  wire  right = _io_redirect_valid_T & ~predictWrong; // @[src/main/scala/nutcore/backend/fu/ALU.scala 176:32]
  wire  _T_55 = right & isBranch; // @[src/main/scala/nutcore/backend/fu/ALU.scala 178:33]
  wire  _T_56 = _io_redirect_valid_T_1 & isBranch; // @[src/main/scala/nutcore/backend/fu/ALU.scala 179:33]
  wire  _T_60 = _T_56 & io_cfIn_pc[2:0] == 3'h0; // @[src/main/scala/nutcore/backend/fu/ALU.scala 180:45]
  wire  _T_61 = _T_56 & io_cfIn_pc[2:0] == 3'h0 & isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 180:73]
  wire  _T_67 = _T_60 & _T_12; // @[src/main/scala/nutcore/backend/fu/ALU.scala 181:73]
  wire  _T_71 = _T_56 & io_cfIn_pc[2:0] == 3'h2; // @[src/main/scala/nutcore/backend/fu/ALU.scala 182:45]
  wire  _T_72 = _T_56 & io_cfIn_pc[2:0] == 3'h2 & isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 182:73]
  wire  _T_78 = _T_71 & _T_12; // @[src/main/scala/nutcore/backend/fu/ALU.scala 183:73]
  wire  _T_82 = _T_56 & io_cfIn_pc[2:0] == 3'h4; // @[src/main/scala/nutcore/backend/fu/ALU.scala 184:45]
  wire  _T_83 = _T_56 & io_cfIn_pc[2:0] == 3'h4 & isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 184:73]
  wire  _T_89 = _T_82 & _T_12; // @[src/main/scala/nutcore/backend/fu/ALU.scala 185:73]
  wire  _T_93 = _T_56 & io_cfIn_pc[2:0] == 3'h6; // @[src/main/scala/nutcore/backend/fu/ALU.scala 186:45]
  wire  _T_94 = _T_56 & io_cfIn_pc[2:0] == 3'h6 & isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 186:73]
  wire  _T_100 = _T_93 & _T_12; // @[src/main/scala/nutcore/backend/fu/ALU.scala 187:73]
  wire  _T_104 = right & _T_21; // @[src/main/scala/nutcore/backend/fu/ALU.scala 188:33]
  wire  _T_108 = _io_redirect_valid_T_1 & _T_21; // @[src/main/scala/nutcore/backend/fu/ALU.scala 189:33]
  wire  _T_110 = right & _T_22; // @[src/main/scala/nutcore/backend/fu/ALU.scala 190:33]
  wire  _T_112 = _io_redirect_valid_T_1 & _T_22; // @[src/main/scala/nutcore/backend/fu/ALU.scala 191:33]
  wire  _T_114 = right & _T_23; // @[src/main/scala/nutcore/backend/fu/ALU.scala 192:33]
  wire  _T_116 = _io_redirect_valid_T_1 & _T_23; // @[src/main/scala/nutcore/backend/fu/ALU.scala 193:33]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  hasIllegalJumpAddr_p; // @[src/main/scala/nutcore/backend/fu/ALU.scala 138:35]
  wire  hasIllegalJumpAddr_t = hasIllegalJumpAddr ^ hasIllegalJumpAddr_p; // @[src/main/scala/nutcore/backend/fu/ALU.scala 138:35]
  wire  toggle_2584_clock;
  wire  toggle_2584_reset;
  wire  toggle_2584_valid;
  reg  toggle_2584_valid_reg;
  reg [63:0] io_jumpIsIllegal_bits_r_p; // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
  wire [63:0] io_jumpIsIllegal_bits_r_t = io_jumpIsIllegal_bits_r ^ io_jumpIsIllegal_bits_r_p; // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
  wire  toggle_2585_clock;
  wire  toggle_2585_reset;
  wire [63:0] toggle_2585_valid;
  reg [63:0] toggle_2585_valid_reg;
  reg  REG_valid_p; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  wire  REG_valid_t = REG_valid ^ REG_valid_p; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  wire  toggle_2649_clock;
  wire  toggle_2649_reset;
  wire  toggle_2649_valid;
  reg  toggle_2649_valid_reg;
  reg [38:0] REG_pc_p; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  wire [38:0] REG_pc_t = REG_pc ^ REG_pc_p; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  wire  toggle_2650_clock;
  wire  toggle_2650_reset;
  wire [38:0] toggle_2650_valid;
  reg [38:0] toggle_2650_valid_reg;
  reg  REG_isMissPredict_p; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  wire  REG_isMissPredict_t = REG_isMissPredict ^ REG_isMissPredict_p; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  wire  toggle_2689_clock;
  wire  toggle_2689_reset;
  wire  toggle_2689_valid;
  reg  toggle_2689_valid_reg;
  reg [38:0] REG_actualTarget_p; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  wire [38:0] REG_actualTarget_t = REG_actualTarget ^ REG_actualTarget_p; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  wire  toggle_2690_clock;
  wire  toggle_2690_reset;
  wire [38:0] toggle_2690_valid;
  reg [38:0] toggle_2690_valid_reg;
  reg  REG_actualTaken_p; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  wire  REG_actualTaken_t = REG_actualTaken ^ REG_actualTaken_p; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  wire  toggle_2729_clock;
  wire  toggle_2729_reset;
  wire  toggle_2729_valid;
  reg  toggle_2729_valid_reg;
  reg [6:0] REG_fuOpType_p; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  wire [6:0] REG_fuOpType_t = REG_fuOpType ^ REG_fuOpType_p; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  wire  toggle_2730_clock;
  wire  toggle_2730_reset;
  wire [6:0] toggle_2730_valid;
  reg [6:0] toggle_2730_valid_reg;
  reg [1:0] REG_btbType_p; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  wire [1:0] REG_btbType_t = REG_btbType ^ REG_btbType_p; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  wire  toggle_2737_clock;
  wire  toggle_2737_reset;
  wire [1:0] toggle_2737_valid;
  reg [1:0] toggle_2737_valid_reg;
  reg  REG_isRVC_p; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  wire  REG_isRVC_t = REG_isRVC ^ REG_isRVC_p; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
  wire  toggle_2739_clock;
  wire  toggle_2739_reset;
  wire  toggle_2739_valid;
  reg  toggle_2739_valid_reg;
  GEN_w1_toggle #(.COVER_INDEX(2584)) toggle_2584 (
    .clock(toggle_2584_clock),
    .reset(toggle_2584_reset),
    .valid(toggle_2584_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(2585)) toggle_2585 (
    .clock(toggle_2585_clock),
    .reset(toggle_2585_reset),
    .valid(toggle_2585_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(2649)) toggle_2649 (
    .clock(toggle_2649_clock),
    .reset(toggle_2649_reset),
    .valid(toggle_2649_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(2650)) toggle_2650 (
    .clock(toggle_2650_clock),
    .reset(toggle_2650_reset),
    .valid(toggle_2650_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(2689)) toggle_2689 (
    .clock(toggle_2689_clock),
    .reset(toggle_2689_reset),
    .valid(toggle_2689_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(2690)) toggle_2690 (
    .clock(toggle_2690_clock),
    .reset(toggle_2690_reset),
    .valid(toggle_2690_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(2729)) toggle_2729 (
    .clock(toggle_2729_clock),
    .reset(toggle_2729_reset),
    .valid(toggle_2729_valid)
  );
  GEN_w7_toggle #(.COVER_INDEX(2730)) toggle_2730 (
    .clock(toggle_2730_clock),
    .reset(toggle_2730_reset),
    .valid(toggle_2730_valid)
  );
  GEN_w2_toggle #(.COVER_INDEX(2737)) toggle_2737 (
    .clock(toggle_2737_clock),
    .reset(toggle_2737_reset),
    .valid(toggle_2737_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(2739)) toggle_2739 (
    .clock(toggle_2739_clock),
    .reset(toggle_2739_reset),
    .valid(toggle_2739_valid)
  );
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/backend/fu/ALU.scala 161:16]
  assign io_out_bits = _io_out_bits_T_10[63:0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 134:15]
  assign io_redirect_target = _io_redirect_target_T_7[38:0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 126:22]
  assign io_redirect_valid = io_in_valid & isBru & predictWrong; // @[src/main/scala/nutcore/backend/fu/ALU.scala 128:39]
  assign io_jumpIsIllegal_valid = hasIllegalJumpAddr; // @[src/main/scala/nutcore/backend/fu/ALU.scala 146:26]
  assign io_jumpIsIllegal_bits = io_jumpIsIllegal_bits_r; // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:25]
  assign REG_0_valid = REG_valid;
  assign REG_0_pc = REG_pc;
  assign REG_0_isMissPredict = REG_isMissPredict;
  assign REG_0_actualTarget = REG_actualTarget;
  assign REG_0_fuOpType = REG_fuOpType;
  assign REG_0_btbType = REG_btbType;
  assign REG_0_isRVC = REG_isRVC;
  assign toggle_2584_clock = clock;
  assign toggle_2584_reset = reset;
  assign toggle_2584_valid = hasIllegalJumpAddr ^ toggle_2584_valid_reg;
  assign toggle_2585_clock = clock;
  assign toggle_2585_reset = reset;
  assign toggle_2585_valid = io_jumpIsIllegal_bits_r ^ toggle_2585_valid_reg;
  assign toggle_2649_clock = clock;
  assign toggle_2649_reset = reset;
  assign toggle_2649_valid = REG_valid ^ toggle_2649_valid_reg;
  assign toggle_2650_clock = clock;
  assign toggle_2650_reset = reset;
  assign toggle_2650_valid = REG_pc ^ toggle_2650_valid_reg;
  assign toggle_2689_clock = clock;
  assign toggle_2689_reset = reset;
  assign toggle_2689_valid = REG_isMissPredict ^ toggle_2689_valid_reg;
  assign toggle_2690_clock = clock;
  assign toggle_2690_reset = reset;
  assign toggle_2690_valid = REG_actualTarget ^ toggle_2690_valid_reg;
  assign toggle_2729_clock = clock;
  assign toggle_2729_reset = reset;
  assign toggle_2729_valid = REG_actualTaken ^ toggle_2729_valid_reg;
  assign toggle_2730_clock = clock;
  assign toggle_2730_reset = reset;
  assign toggle_2730_valid = REG_fuOpType ^ toggle_2730_valid_reg;
  assign toggle_2737_clock = clock;
  assign toggle_2737_reset = reset;
  assign toggle_2737_valid = REG_btbType ^ toggle_2737_valid_reg;
  assign toggle_2739_clock = clock;
  assign toggle_2739_reset = reset;
  assign toggle_2739_valid = REG_isRVC ^ toggle_2739_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/ALU.scala 138:35]
      hasIllegalJumpAddr <= 1'h0; // @[src/main/scala/nutcore/backend/fu/ALU.scala 138:35]
    end else begin
      hasIllegalJumpAddr <= _GEN_1;
    end
    if (isIllegalJumpAddr) begin // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
      if (isBranch) begin // @[src/main/scala/nutcore/backend/fu/ALU.scala 121:19]
        io_jumpIsIllegal_bits_r <= _target_T_3;
      end else begin
        io_jumpIsIllegal_bits_r <= _target_T_5;
      end
    end
    REG_valid <= io_in_valid & isBru; // @[src/main/scala/nutcore/backend/fu/ALU.scala 164:31]
    REG_pc <= io_cfIn_pc; // @[src/main/scala/nutcore/backend/fu/ALU.scala 163:30 165:19]
    if (~taken & isBranch) begin // @[src/main/scala/nutcore/backend/fu/ALU.scala 122:25]
      REG_isMissPredict <= io_cfIn_brIdx[0];
    end else begin
      REG_isMissPredict <= ~io_cfIn_brIdx[0] | io_redirect_target != io_cfIn_pnpc;
    end
    REG_actualTarget <= target[38:0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 163:30 167:29]
    REG_actualTaken <= _taken_T_8 ^ io_in_bits_func[0]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 120:72]
    REG_fuOpType <= io_in_bits_func; // @[src/main/scala/nutcore/backend/fu/ALU.scala 163:30 169:25]
    REG_btbType <= _T_53 | _T_45; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
    REG_isRVC <= io_cfIn_instr[1:0] != 2'h3; // @[src/main/scala/nutcore/backend/fu/ALU.scala 123:35]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_cfIn_instr[1:0] == 2'h3 | isRVC | ~io_in_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ALU.scala:124 assert(io.cfIn.instr(1,0) === \"b11\".U || isRVC || !valid)\n"); // @[src/main/scala/nutcore/backend/fu/ALU.scala 124:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    hasIllegalJumpAddr_p <= hasIllegalJumpAddr; // @[src/main/scala/nutcore/backend/fu/ALU.scala 138:35]
    toggle_2584_valid_reg <= hasIllegalJumpAddr;
    io_jumpIsIllegal_bits_r_p <= io_jumpIsIllegal_bits_r; // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    toggle_2585_valid_reg <= io_jumpIsIllegal_bits_r;
    REG_valid_p <= REG_valid; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    toggle_2649_valid_reg <= REG_valid;
    REG_pc_p <= REG_pc; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    toggle_2650_valid_reg <= REG_pc;
    REG_isMissPredict_p <= REG_isMissPredict; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    toggle_2689_valid_reg <= REG_isMissPredict;
    REG_actualTarget_p <= REG_actualTarget; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    toggle_2690_valid_reg <= REG_actualTarget;
    REG_actualTaken_p <= REG_actualTaken; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    toggle_2729_valid_reg <= REG_actualTaken;
    REG_fuOpType_p <= REG_fuOpType; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    toggle_2730_valid_reg <= REG_fuOpType;
    REG_btbType_p <= REG_btbType; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    toggle_2737_valid_reg <= REG_btbType;
    REG_isRVC_p <= REG_isRVC; // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    toggle_2739_valid_reg <= REG_isRVC;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  hasIllegalJumpAddr = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  io_jumpIsIllegal_bits_r = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  REG_valid = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  REG_pc = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  REG_isMissPredict = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  REG_actualTarget = _RAND_5[38:0];
  _RAND_6 = {1{`RANDOM}};
  REG_actualTaken = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  REG_fuOpType = _RAND_7[6:0];
  _RAND_8 = {1{`RANDOM}};
  REG_btbType = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  REG_isRVC = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  hasIllegalJumpAddr_p = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  toggle_2584_valid_reg = _RAND_11[0:0];
  _RAND_12 = {2{`RANDOM}};
  io_jumpIsIllegal_bits_r_p = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  toggle_2585_valid_reg = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  REG_valid_p = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  toggle_2649_valid_reg = _RAND_15[0:0];
  _RAND_16 = {2{`RANDOM}};
  REG_pc_p = _RAND_16[38:0];
  _RAND_17 = {2{`RANDOM}};
  toggle_2650_valid_reg = _RAND_17[38:0];
  _RAND_18 = {1{`RANDOM}};
  REG_isMissPredict_p = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  toggle_2689_valid_reg = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  REG_actualTarget_p = _RAND_20[38:0];
  _RAND_21 = {2{`RANDOM}};
  toggle_2690_valid_reg = _RAND_21[38:0];
  _RAND_22 = {1{`RANDOM}};
  REG_actualTaken_p = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  toggle_2729_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  REG_fuOpType_p = _RAND_24[6:0];
  _RAND_25 = {1{`RANDOM}};
  toggle_2730_valid_reg = _RAND_25[6:0];
  _RAND_26 = {1{`RANDOM}};
  REG_btbType_p = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  toggle_2737_valid_reg = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  REG_isRVC_p = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  toggle_2739_valid_reg = _RAND_29[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(io_cfIn_instr[1:0] == 2'h3 | isRVC | ~io_in_valid); // @[src/main/scala/nutcore/backend/fu/ALU.scala 124:9]
    end
    //
    if (enToggle_past) begin
      cover(hasIllegalJumpAddr_t); // @[src/main/scala/nutcore/backend/fu/ALU.scala 138:35]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[0]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[1]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[2]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[3]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[4]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[5]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[6]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[7]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[8]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[9]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[10]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[11]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[12]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[13]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[14]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[15]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[16]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[17]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[18]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[19]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[20]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[21]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[22]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[23]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[24]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[25]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[26]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[27]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[28]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[29]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[30]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[31]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[32]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[33]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[34]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[35]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[36]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[37]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[38]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[39]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[40]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[41]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[42]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[43]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[44]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[45]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[46]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[47]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[48]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[49]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[50]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[51]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[52]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[53]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[54]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[55]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[56]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[57]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[58]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[59]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[60]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[61]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[62]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(io_jumpIsIllegal_bits_r_t[63]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 147:37]
    end
    //
    if (enToggle_past) begin
      cover(REG_valid_t); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[0]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[1]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[2]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[3]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[4]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[5]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[6]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[7]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[8]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[9]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[10]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[11]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[12]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[13]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[14]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[15]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[16]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[17]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[18]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[19]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[20]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[21]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[22]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[23]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[24]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[25]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[26]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[27]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[28]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[29]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[30]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[31]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[32]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[33]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[34]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[35]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[36]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[37]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_pc_t[38]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_isMissPredict_t); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[0]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[1]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[2]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[3]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[4]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[5]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[6]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[7]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[8]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[9]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[10]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[11]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[12]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[13]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[14]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[15]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[16]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[17]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[18]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[19]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[20]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[21]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[22]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[23]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[24]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[25]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[26]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[27]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[28]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[29]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[30]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[31]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[32]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[33]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[34]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[35]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[36]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[37]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTarget_t[38]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_actualTaken_t); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_fuOpType_t[0]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_fuOpType_t[1]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_fuOpType_t[2]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_fuOpType_t[3]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_fuOpType_t[4]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_fuOpType_t[5]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_fuOpType_t[6]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_btbType_t[0]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_btbType_t[1]); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
    //
    if (enToggle_past) begin
      cover(REG_isRVC_t); // @[src/main/scala/nutcore/backend/fu/ALU.scala 174:34]
    end
  end
endmodule
module LSExecUnit(
  input         clock,
  input         reset,
  output        io__in_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input         io__in_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input  [63:0] io__in_bits_src1, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input  [6:0]  io__in_bits_func, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input         io__out_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__out_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [63:0] io__out_bits, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input  [63:0] io__wdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input         io__dmem_req_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__dmem_req_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [38:0] io__dmem_req_bits_addr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [2:0]  io__dmem_req_bits_size, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [3:0]  io__dmem_req_bits_cmd, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [7:0]  io__dmem_req_bits_wmask, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [63:0] io__dmem_req_bits_wdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__dmem_resp_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input         io__dmem_resp_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input  [63:0] io__dmem_resp_bits_rdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__isMMIO, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__dtlbPF, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__dtlbAF, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output [63:0] io__vaddr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__loadAccessFault, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  output        io__storeAccessFault, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 377:14]
  input         DTLBPF,
  input         scIsSuccess_0,
  input         vmEnable_0,
  input         ISAMO2,
  input         DTLBFINISH,
  input         DTLBAF
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  _io_vaddr_T = io__in_ready & io__in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg [63:0] io_vaddr_r; // @[src/main/scala/utils/Hold.scala 23:65]
  reg [63:0] addrLatch; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
  wire  isStore = io__in_valid & io__in_bits_func[3]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 423:23]
  wire  partialLoad = ~isStore & io__in_bits_func != 7'h3; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 424:30]
  reg [1:0] state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 427:22]
  wire [5:0] vaddrPF_lo_lo = {io__vaddr[58] != io__vaddr[38],io__vaddr[59] != io__vaddr[38],io__vaddr[60] != io__vaddr[
    38],io__vaddr[61] != io__vaddr[38],io__vaddr[62] != io__vaddr[38],io__vaddr[63] != io__vaddr[38]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 442:43]
  wire [11:0] vaddrPF_lo = {io__vaddr[52] != io__vaddr[38],io__vaddr[53] != io__vaddr[38],io__vaddr[54] != io__vaddr[38]
    ,io__vaddr[55] != io__vaddr[38],io__vaddr[56] != io__vaddr[38],io__vaddr[57] != io__vaddr[38],vaddrPF_lo_lo}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 442:43]
  wire [5:0] vaddrPF_hi_lo = {io__vaddr[46] != io__vaddr[38],io__vaddr[47] != io__vaddr[38],io__vaddr[48] != io__vaddr[
    38],io__vaddr[49] != io__vaddr[38],io__vaddr[50] != io__vaddr[38],io__vaddr[51] != io__vaddr[38]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 442:43]
  wire [24:0] _vaddrPF_T_76 = {io__vaddr[39] != io__vaddr[38],io__vaddr[40] != io__vaddr[38],io__vaddr[41] != io__vaddr[
    38],io__vaddr[42] != io__vaddr[38],io__vaddr[43] != io__vaddr[38],io__vaddr[44] != io__vaddr[38],io__vaddr[45] !=
    io__vaddr[38],vaddrPF_hi_lo,vaddrPF_lo}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 442:43]
  wire  vaddrPF = io__in_valid & vmEnable_0 & |_vaddrPF_T_76; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 442:37]
  wire  dtlbHasException = DTLBPF | DTLBAF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 446:33]
  wire  _T_1 = io__dmem_req_ready & io__dmem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_4 = ~vmEnable_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 450:32]
  wire [1:0] _GEN_3 = DTLBFINISH & (dtlbHasException | ~scIsSuccess_0) ? 2'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 427:22 454:{63,71}]
  wire  _T_14 = io__dmem_resp_ready & io__dmem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [1:0] _state_T = partialLoad ? 2'h3 : 2'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 457:62]
  wire [1:0] _GEN_5 = _T_14 ? _state_T : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 427:22 457:{48,56}]
  wire [1:0] _GEN_6 = 2'h3 == state ? 2'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 447:18 427:22 458:32]
  wire [63:0] _reqWdata_T_3 = {io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0]
    ,io__wdata[7:0],io__wdata[7:0]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 399:22]
  wire [63:0] _reqWdata_T_6 = {io__wdata[15:0],io__wdata[15:0],io__wdata[15:0],io__wdata[15:0]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 400:22]
  wire [63:0] _reqWdata_T_8 = {io__wdata[31:0],io__wdata[31:0]}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 401:22]
  wire  _reqWdata_T_9 = 2'h0 == io__in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _reqWdata_T_10 = 2'h1 == io__in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _reqWdata_T_11 = 2'h2 == io__in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _reqWdata_T_12 = 2'h3 == io__in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _reqWdata_T_13 = _reqWdata_T_9 ? _reqWdata_T_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_14 = _reqWdata_T_10 ? _reqWdata_T_6 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_15 = _reqWdata_T_11 ? _reqWdata_T_8 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_16 = _reqWdata_T_12 ? io__wdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_17 = _reqWdata_T_13 | _reqWdata_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _reqWdata_T_18 = _reqWdata_T_17 | _reqWdata_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _reqWmask_T_5 = _reqWdata_T_10 ? 2'h3 : 2'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _reqWmask_T_6 = _reqWdata_T_11 ? 4'hf : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _reqWmask_T_7 = _reqWdata_T_12 ? 8'hff : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _GEN_20 = {{1'd0}, _reqWdata_T_9}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [1:0] _reqWmask_T_8 = _GEN_20 | _reqWmask_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _GEN_21 = {{2'd0}, _reqWmask_T_8}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _reqWmask_T_9 = _GEN_21 | _reqWmask_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _GEN_22 = {{4'd0}, _reqWmask_T_9}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _reqWmask_T_10 = _GEN_22 | _reqWmask_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [14:0] _GEN_30 = {{7'd0}, _reqWmask_T_10}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 395:8]
  wire [14:0] reqWmask = _GEN_30 << io__in_bits_src1[2:0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 395:8]
  wire  hasException = io__loadAccessFault | io__storeAccessFault | vaddrPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 476:64]
  wire  _io_dmem_req_valid_T = state == 2'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 477:37]
  wire  _io_out_valid_T_3 = state == 2'h3; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 483:13]
  wire  _io_out_valid_T_6 = _T_14 & state == 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 484:22]
  wire  _io_out_valid_T_7 = partialLoad ? _io_out_valid_T_3 : _io_out_valid_T_6; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 482:8]
  reg [63:0] rdataLatch; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
  wire  _rdataSel64_T_9 = 3'h0 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_10 = 3'h1 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_11 = 3'h2 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_12 = 3'h3 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_13 = 3'h4 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_14 = 3'h5 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_15 = 3'h6 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataSel64_T_16 = 3'h7 == addrLatch[2:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdataSel64_T_17 = _rdataSel64_T_9 ? rdataLatch : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [55:0] _rdataSel64_T_18 = _rdataSel64_T_10 ? rdataLatch[63:8] : 56'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [47:0] _rdataSel64_T_19 = _rdataSel64_T_11 ? rdataLatch[63:16] : 48'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [39:0] _rdataSel64_T_20 = _rdataSel64_T_12 ? rdataLatch[63:24] : 40'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdataSel64_T_21 = _rdataSel64_T_13 ? rdataLatch[63:32] : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [23:0] _rdataSel64_T_22 = _rdataSel64_T_14 ? rdataLatch[63:40] : 24'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [15:0] _rdataSel64_T_23 = _rdataSel64_T_15 ? rdataLatch[63:48] : 16'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _rdataSel64_T_24 = _rdataSel64_T_16 ? rdataLatch[63:56] : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_23 = {{8'd0}, _rdataSel64_T_18}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_25 = _rdataSel64_T_17 | _GEN_23; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_24 = {{16'd0}, _rdataSel64_T_19}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_26 = _rdataSel64_T_25 | _GEN_24; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_25 = {{24'd0}, _rdataSel64_T_20}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_27 = _rdataSel64_T_26 | _GEN_25; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_26 = {{32'd0}, _rdataSel64_T_21}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_28 = _rdataSel64_T_27 | _GEN_26; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_27 = {{40'd0}, _rdataSel64_T_22}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_29 = _rdataSel64_T_28 | _GEN_27; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_28 = {{48'd0}, _rdataSel64_T_23}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataSel64_T_30 = _rdataSel64_T_29 | _GEN_28; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _GEN_29 = {{56'd0}, _rdataSel64_T_24}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdataSel64 = _rdataSel64_T_30 | _GEN_29; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  rdataPartialLoad_signBit = rdataSel64[7]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [55:0] _rdataPartialLoad_T_1 = rdataPartialLoad_signBit ? 56'hffffffffffffff : 56'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _rdataPartialLoad_T_2 = {_rdataPartialLoad_T_1,rdataSel64[7:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  rdataPartialLoad_signBit_1 = rdataSel64[15]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [47:0] _rdataPartialLoad_T_4 = rdataPartialLoad_signBit_1 ? 48'hffffffffffff : 48'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _rdataPartialLoad_T_5 = {_rdataPartialLoad_T_4,rdataSel64[15:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  rdataPartialLoad_signBit_2 = rdataSel64[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _rdataPartialLoad_T_7 = rdataPartialLoad_signBit_2 ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _rdataPartialLoad_T_8 = {_rdataPartialLoad_T_7,rdataSel64[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _rdataPartialLoad_T_10 = {56'h0,rdataSel64[7:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _rdataPartialLoad_T_12 = {48'h0,rdataSel64[15:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _rdataPartialLoad_T_14 = {32'h0,rdataSel64[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  _rdataPartialLoad_T_15 = 7'h0 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_16 = 7'h1 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_17 = 7'h2 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_18 = 7'h4 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_19 = 7'h5 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdataPartialLoad_T_20 = 7'h6 == io__in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdataPartialLoad_T_21 = _rdataPartialLoad_T_15 ? _rdataPartialLoad_T_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_22 = _rdataPartialLoad_T_16 ? _rdataPartialLoad_T_5 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_23 = _rdataPartialLoad_T_17 ? _rdataPartialLoad_T_8 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_24 = _rdataPartialLoad_T_18 ? _rdataPartialLoad_T_10 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_25 = _rdataPartialLoad_T_19 ? _rdataPartialLoad_T_12 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_26 = _rdataPartialLoad_T_20 ? _rdataPartialLoad_T_14 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_27 = _rdataPartialLoad_T_21 | _rdataPartialLoad_T_22; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_28 = _rdataPartialLoad_T_27 | _rdataPartialLoad_T_23; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_29 = _rdataPartialLoad_T_28 | _rdataPartialLoad_T_24; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdataPartialLoad_T_30 = _rdataPartialLoad_T_29 | _rdataPartialLoad_T_25; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdataPartialLoad = _rdataPartialLoad_T_30 | _rdataPartialLoad_T_26; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_loadAccessFault_T_1 = io__in_valid & _T_4; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 531:32]
  wire  _io_loadAccessFault_T_7 = io__in_bits_src1 >= 64'h38000000 & io__in_bits_src1 < 64'h38010000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_10 = io__in_bits_src1 >= 64'h3c000000 & io__in_bits_src1 < 64'h40000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_13 = io__in_bits_src1 >= 64'h40600000 & io__in_bits_src1 < 64'h40600010; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_16 = io__in_bits_src1 >= 64'h50000000 & io__in_bits_src1 < 64'h50400000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_19 = io__in_bits_src1 >= 64'h40001000 & io__in_bits_src1 < 64'h40001008; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_22 = io__in_bits_src1 >= 64'h40000000 & io__in_bits_src1 < 64'h40001000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_25 = io__in_bits_src1 >= 64'h40002000 & io__in_bits_src1 < 64'h40003000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _io_loadAccessFault_T_28 = io__in_bits_src1 >= 64'h80000000 & io__in_bits_src1 < 64'h100000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [7:0] _io_loadAccessFault_T_29 = {_io_loadAccessFault_T_28,_io_loadAccessFault_T_25,_io_loadAccessFault_T_22,
    _io_loadAccessFault_T_19,_io_loadAccessFault_T_16,_io_loadAccessFault_T_13,_io_loadAccessFault_T_10,
    _io_loadAccessFault_T_7}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _io_loadAccessFault_T_30 = |_io_loadAccessFault_T_29; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  _io_loadAccessFault_T_31 = ~_io_loadAccessFault_T_30; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 531:71]
  wire  _io_storeAccessFault_T_33 = |(io__in_bits_src1 >= 64'h80000000 & io__in_bits_src1 < 64'h100000000); // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  _T_30 = ~io__dmem_req_bits_cmd[0] & ~io__dmem_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _T_31 = io__dmem_req_valid & _T_30; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  wire  _T_33 = _T_31 & _T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 534:39]
  reg  r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_10 = _T_31 | r; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _T_42 = io__dmem_req_valid & io__dmem_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  reg  r_1; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_12 = _T_42 | r_1; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [63:0] io_vaddr_r_p; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [63:0] io_vaddr_r_t = io_vaddr_r ^ io_vaddr_r_p; // @[src/main/scala/utils/Hold.scala 23:65]
  wire  toggle_2740_clock;
  wire  toggle_2740_reset;
  wire [63:0] toggle_2740_valid;
  reg [63:0] toggle_2740_valid_reg;
  reg [63:0] addrLatch_p; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
  wire [63:0] addrLatch_t = addrLatch ^ addrLatch_p; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
  wire  toggle_2804_clock;
  wire  toggle_2804_reset;
  wire [63:0] toggle_2804_valid;
  reg [63:0] toggle_2804_valid_reg;
  reg [1:0] state_p; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 427:22]
  wire [1:0] state_t = state ^ state_p; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 427:22]
  wire  toggle_2868_clock;
  wire  toggle_2868_reset;
  wire [1:0] toggle_2868_valid;
  reg [1:0] toggle_2868_valid_reg;
  reg [63:0] rdataLatch_p; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
  wire [63:0] rdataLatch_t = rdataLatch ^ rdataLatch_p; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
  wire  toggle_2870_clock;
  wire  toggle_2870_reset;
  wire [63:0] toggle_2870_valid;
  reg [63:0] toggle_2870_valid_reg;
  reg  r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  r_t = r ^ r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_2934_clock;
  wire  toggle_2934_reset;
  wire  toggle_2934_valid;
  reg  toggle_2934_valid_reg;
  reg  r_1_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  r_1_t = r_1 ^ r_1_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_2935_clock;
  wire  toggle_2935_reset;
  wire  toggle_2935_valid;
  reg  toggle_2935_valid_reg;
  GEN_w64_toggle #(.COVER_INDEX(2740)) toggle_2740 (
    .clock(toggle_2740_clock),
    .reset(toggle_2740_reset),
    .valid(toggle_2740_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(2804)) toggle_2804 (
    .clock(toggle_2804_clock),
    .reset(toggle_2804_reset),
    .valid(toggle_2804_valid)
  );
  GEN_w2_toggle #(.COVER_INDEX(2868)) toggle_2868 (
    .clock(toggle_2868_clock),
    .reset(toggle_2868_reset),
    .valid(toggle_2868_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(2870)) toggle_2870 (
    .clock(toggle_2870_clock),
    .reset(toggle_2870_reset),
    .valid(toggle_2870_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(2934)) toggle_2934 (
    .clock(toggle_2934_clock),
    .reset(toggle_2934_reset),
    .valid(toggle_2934_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(2935)) toggle_2935 (
    .clock(toggle_2935_clock),
    .reset(toggle_2935_reset),
    .valid(toggle_2935_valid)
  );
  assign io__in_ready = _io_dmem_req_valid_T | dtlbHasException; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 487:37]
  assign io__out_valid = dtlbHasException & state != 2'h0 | hasException | _io_out_valid_T_7; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 480:22]
  assign io__out_bits = partialLoad ? rdataPartialLoad : io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 520:21]
  assign io__dmem_req_valid = io__in_valid & state == 2'h0 & ~hasException; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 477:49]
  assign io__dmem_req_bits_addr = io__in_bits_src1[38:0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 466:68]
  assign io__dmem_req_bits_size = {{1'd0}, io__in_bits_func[1:0]}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 66:15]
  assign io__dmem_req_bits_cmd = {{3'd0}, isStore}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io__dmem_req_bits_wmask = reqWmask[7:0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 68:16]
  assign io__dmem_req_bits_wdata = _reqWdata_T_18 | _reqWdata_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io__dmem_resp_ready = 1'h1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 478:19]
  assign io__isMMIO = 1'h0;
  assign io__dtlbPF = DTLBPF | vaddrPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 443:23]
  assign io__dtlbAF = DTLBAF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 431:24]
  assign io__vaddr = _io_vaddr_T ? io__in_bits_src1 : io_vaddr_r; // @[src/main/scala/utils/Hold.scala 23:48]
  assign io__loadAccessFault = io__in_valid & _T_4 & ~(isStore | ISAMO2) & ~_io_loadAccessFault_T_30; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 531:68]
  assign io__storeAccessFault = _io_loadAccessFault_T_1 & (isStore & _io_loadAccessFault_T_31 | ISAMO2 & ~
    _io_storeAccessFault_T_33); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 532:45]
  assign toggle_2740_clock = clock;
  assign toggle_2740_reset = reset;
  assign toggle_2740_valid = io_vaddr_r ^ toggle_2740_valid_reg;
  assign toggle_2804_clock = clock;
  assign toggle_2804_reset = reset;
  assign toggle_2804_valid = addrLatch ^ toggle_2804_valid_reg;
  assign toggle_2868_clock = clock;
  assign toggle_2868_reset = reset;
  assign toggle_2868_valid = state ^ toggle_2868_valid_reg;
  assign toggle_2870_clock = clock;
  assign toggle_2870_reset = reset;
  assign toggle_2870_valid = rdataLatch ^ toggle_2870_valid_reg;
  assign toggle_2934_clock = clock;
  assign toggle_2934_reset = reset;
  assign toggle_2934_valid = r ^ toggle_2934_valid_reg;
  assign toggle_2935_clock = clock;
  assign toggle_2935_reset = reset;
  assign toggle_2935_valid = r_1 ^ toggle_2935_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      io_vaddr_r <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_io_vaddr_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      io_vaddr_r <= io__in_bits_src1; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    addrLatch <= io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 427:22]
      state <= 2'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 427:22]
    end else if (2'h0 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 447:18]
      if (_T_1 & ~vmEnable_0) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 450:45]
        state <= 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 450:53]
      end else if (_T_1 & vmEnable_0) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 449:45]
        state <= 2'h1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 449:53]
      end
    end else if (2'h1 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 447:18]
      if (DTLBFINISH & ~dtlbHasException & scIsSuccess_0) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 455:61]
        state <= 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 455:69]
      end else begin
        state <= _GEN_3;
      end
    end else if (2'h2 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 447:18]
      state <= _GEN_5;
    end else begin
      state <= _GEN_6;
    end
    rdataLatch <= io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (_T_14) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      r <= _GEN_10;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_1 <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (_T_14) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      r_1 <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      r_1 <= _GEN_12;
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    io_vaddr_r_p <= io_vaddr_r; // @[src/main/scala/utils/Hold.scala 23:65]
    toggle_2740_valid_reg <= io_vaddr_r;
    addrLatch_p <= addrLatch; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    toggle_2804_valid_reg <= addrLatch;
    state_p <= state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 427:22]
    toggle_2868_valid_reg <= state;
    rdataLatch_p <= rdataLatch; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    toggle_2870_valid_reg <= rdataLatch;
    r_p <= r; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_2934_valid_reg <= r;
    r_1_p <= r_1; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_2935_valid_reg <= r_1;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  io_vaddr_r = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  addrLatch = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[1:0];
  _RAND_3 = {2{`RANDOM}};
  rdataLatch = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  r_1 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  io_vaddr_r_p = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  toggle_2740_valid_reg = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  addrLatch_p = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  toggle_2804_valid_reg = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  state_p = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  toggle_2868_valid_reg = _RAND_11[1:0];
  _RAND_12 = {2{`RANDOM}};
  rdataLatch_p = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  toggle_2870_valid_reg = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  r_p = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  toggle_2934_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  r_1_p = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  toggle_2935_valid_reg = _RAND_17[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[0]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[1]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[2]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[3]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[4]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[5]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[6]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[7]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[8]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[9]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[10]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[11]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[12]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[13]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[14]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[15]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[16]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[17]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[18]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[19]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[20]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[21]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[22]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[23]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[24]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[25]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[26]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[27]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[28]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[29]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[30]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[31]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[32]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[33]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[34]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[35]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[36]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[37]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[38]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[39]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[40]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[41]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[42]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[43]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[44]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[45]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[46]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[47]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[48]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[49]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[50]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[51]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[52]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[53]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[54]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[55]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[56]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[57]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[58]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[59]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[60]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[61]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[62]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[63]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[0]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[1]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[2]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[3]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[4]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[5]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[6]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[7]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[8]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[9]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[10]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[11]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[12]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[13]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[14]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[15]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[16]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[17]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[18]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[19]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[20]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[21]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[22]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[23]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[24]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[25]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[26]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[27]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[28]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[29]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[30]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[31]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[32]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[33]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[34]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[35]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[36]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[37]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[38]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[39]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[40]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[41]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[42]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[43]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[44]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[45]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[46]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[47]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[48]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[49]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[50]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[51]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[52]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[53]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[54]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[55]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[56]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[57]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[58]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[59]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[60]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[61]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[62]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(addrLatch_t[63]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 422:26]
    end
    //
    if (enToggle_past) begin
      cover(state_t[0]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 427:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[1]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 427:22]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[0]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[1]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[2]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[3]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[4]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[5]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[6]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[7]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[8]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[9]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[10]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[11]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[12]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[13]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[14]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[15]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[16]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[17]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[18]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[19]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[20]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[21]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[22]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[23]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[24]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[25]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[26]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[27]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[28]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[29]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[30]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[31]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[32]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[33]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[34]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[35]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[36]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[37]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[38]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[39]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[40]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[41]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[42]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[43]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[44]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[45]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[46]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[47]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[48]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[49]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[50]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[51]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[52]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[53]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[54]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[55]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[56]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[57]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[58]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[59]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[60]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[61]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[62]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(rdataLatch_t[63]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 492:27]
    end
    //
    if (enToggle_past) begin
      cover(r_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
  end
endmodule
module AtomALU(
  input         clock,
  input         reset,
  input  [63:0] io_src1, // @[src/main/scala/nutcore/backend/fu/LSU.scala 173:14]
  input  [63:0] io_src2, // @[src/main/scala/nutcore/backend/fu/LSU.scala 173:14]
  input  [6:0]  io_func, // @[src/main/scala/nutcore/backend/fu/LSU.scala 173:14]
  input         io_isWordOp, // @[src/main/scala/nutcore/backend/fu/LSU.scala 173:14]
  output [63:0] io_result // @[src/main/scala/nutcore/backend/fu/LSU.scala 173:14]
);
  wire  src1_signBit = io_src1[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _src1_T_1 = src1_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _src1_T_2 = {_src1_T_1,io_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] src1 = io_isWordOp ? _src1_T_2 : io_src1; // @[src/main/scala/nutcore/backend/fu/LSU.scala 183:17]
  wire  src2_signBit = io_src2[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _src2_T_1 = src2_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _src2_T_2 = {_src2_T_1,io_src2[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] src2 = io_isWordOp ? _src2_T_2 : io_src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 184:17]
  wire  isAdderSub = ~io_func[6]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 186:20]
  wire [63:0] _adderRes_T = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[src/main/scala/nutcore/backend/fu/LSU.scala 187:39]
  wire [63:0] _adderRes_T_1 = src2 ^ _adderRes_T; // @[src/main/scala/nutcore/backend/fu/LSU.scala 187:33]
  wire [64:0] _adderRes_T_2 = src1 + _adderRes_T_1; // @[src/main/scala/nutcore/backend/fu/LSU.scala 187:24]
  wire [64:0] _GEN_0 = {{64'd0}, isAdderSub}; // @[src/main/scala/nutcore/backend/fu/LSU.scala 187:60]
  wire [64:0] adderRes = _adderRes_T_2 + _GEN_0; // @[src/main/scala/nutcore/backend/fu/LSU.scala 187:60]
  wire [63:0] xorRes = src1 ^ src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 188:21]
  wire  sltu = ~adderRes[64]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 189:14]
  wire  slt = xorRes[63] ^ sltu; // @[src/main/scala/nutcore/backend/fu/LSU.scala 190:28]
  wire [63:0] _res_T_1 = src1 & src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 196:32]
  wire [63:0] _res_T_2 = src1 | src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 197:32]
  wire [63:0] _res_T_4 = slt ? src1 : src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 198:29]
  wire [63:0] _res_T_6 = slt ? src2 : src1; // @[src/main/scala/nutcore/backend/fu/LSU.scala 199:29]
  wire [63:0] _res_T_8 = sltu ? src1 : src2; // @[src/main/scala/nutcore/backend/fu/LSU.scala 200:29]
  wire [63:0] _res_T_10 = sltu ? src2 : src1; // @[src/main/scala/nutcore/backend/fu/LSU.scala 201:29]
  wire [64:0] _res_T_12 = 6'h22 == io_func[5:0] ? {{1'd0}, src2} : adderRes; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_14 = 6'h24 == io_func[5:0] ? {{1'd0}, xorRes} : _res_T_12; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_16 = 6'h25 == io_func[5:0] ? {{1'd0}, _res_T_1} : _res_T_14; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_18 = 6'h26 == io_func[5:0] ? {{1'd0}, _res_T_2} : _res_T_16; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_20 = 6'h37 == io_func[5:0] ? {{1'd0}, _res_T_4} : _res_T_18; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_22 = 6'h30 == io_func[5:0] ? {{1'd0}, _res_T_6} : _res_T_20; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] _res_T_24 = 6'h31 == io_func[5:0] ? {{1'd0}, _res_T_8} : _res_T_22; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [64:0] res = 6'h32 == io_func[5:0] ? {{1'd0}, _res_T_10} : _res_T_24; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  assign io_result = res[63:0]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 204:13]
endmodule
module UnpipelinedLSU(
  input         clock,
  input         reset,
  input         io__in_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input  [63:0] io__in_bits_src1, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input  [63:0] io__in_bits_src2, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input  [6:0]  io__in_bits_func, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input         io__out_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__out_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [63:0] io__out_bits, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input  [63:0] io__wdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input  [31:0] io__instr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input         io__dmem_req_ready, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__dmem_req_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [38:0] io__dmem_req_bits_addr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [2:0]  io__dmem_req_bits_size, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [3:0]  io__dmem_req_bits_cmd, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [7:0]  io__dmem_req_bits_wmask, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [63:0] io__dmem_req_bits_wdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input         io__dmem_resp_valid, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  input  [63:0] io__dmem_resp_bits_rdata, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__isMMIO, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__dtlbPF, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__dtlbAF, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output [63:0] io__vaddr, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__loadAddrMisaligned, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__storeAddrMisaligned, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__loadAccessFault, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        io__storeAccessFault, // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 45:14]
  output        setLr_0,
  input         lr_0,
  output        scInflight_0,
  output        amoReq_0,
  input  [63:0] lr_addr,
  input  [55:0] dtlb_paddr,
  input         _T_12_0,
  input         scIsSuccess_0,
  output        setLrVal_0,
  input         vmEnable,
  input         DTLBFINISH,
  input         lsuMMIO_0,
  input         _T_13_1,
  output [63:0] setLrAddr_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire  lsExecUnit_clock; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_reset; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__in_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__in_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [63:0] lsExecUnit_io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [6:0] lsExecUnit_io__in_bits_func; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__out_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__out_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [63:0] lsExecUnit_io__out_bits; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [63:0] lsExecUnit_io__wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__dmem_req_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [38:0] lsExecUnit_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [2:0] lsExecUnit_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [3:0] lsExecUnit_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [7:0] lsExecUnit_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [63:0] lsExecUnit_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__dmem_resp_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [63:0] lsExecUnit_io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__isMMIO; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__dtlbPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__dtlbAF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire [63:0] lsExecUnit_io__vaddr; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__loadAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_io__storeAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_DTLBPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_scIsSuccess_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_vmEnable_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_ISAMO2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_DTLBFINISH; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  lsExecUnit_DTLBAF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
  wire  atomALU_clock; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
  wire  atomALU_reset; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
  wire [63:0] atomALU_io_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
  wire [63:0] atomALU_io_src2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
  wire [6:0] atomALU_io_func; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
  wire  atomALU_io_isWordOp; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
  wire [63:0] atomALU_io_result; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
  wire  isAtomic = io__in_bits_func[5]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 54:38]
  wire  _isAmo_T_1 = io__in_bits_func == 7'h20; // @[src/main/scala/nutcore/backend/fu/LSU.scala 57:37]
  wire  _isAmo_T_4 = io__in_bits_func == 7'h21; // @[src/main/scala/nutcore/backend/fu/LSU.scala 58:37]
  wire  isAmo = isAtomic & ~_isAmo_T_1 & ~_isAmo_T_4; // @[src/main/scala/nutcore/backend/fu/LSU.scala 59:61]
  wire [63:0] _in_vaddr_T_1 = io__in_bits_src1 + io__in_bits_src2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 62:43]
  wire [63:0] in_vaddr = isAtomic ? io__in_bits_src1 : _in_vaddr_T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 62:21]
  wire [1:0] _in_func_T_1 = io__instr[12] ? 2'h3 : 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 66:34]
  wire [1:0] in_func = isAtomic ? _in_func_T_1 : io__in_bits_func[1:0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 66:20]
  wire  _addrAligned_T_1 = ~in_vaddr[0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 69:29]
  wire  _addrAligned_T_3 = in_vaddr[1:0] == 2'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 70:32]
  wire  _addrAligned_T_5 = in_vaddr[2:0] == 3'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 71:32]
  wire  _addrAligned_T_6 = 2'h0 == in_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _addrAligned_T_7 = 2'h1 == in_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _addrAligned_T_8 = 2'h2 == in_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _addrAligned_T_9 = 2'h3 == in_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  addrAligned = _addrAligned_T_6 | _addrAligned_T_7 & _addrAligned_T_1 | _addrAligned_T_8 & _addrAligned_T_3 |
    _addrAligned_T_9 & _addrAligned_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  hasAddrMisaligned = io__in_valid & ~addrAligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 73:36]
  wire  _io_loadAddrMisaligned_T_4 = ~io__in_bits_func[3] & ~isAtomic; // @[src/main/scala/nutcore/backend/fu/LSU.scala 56:49]
  wire  _hasScAccessFault_T_1 = ~vmEnable; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 84:46]
  wire  _hasScAccessFault_T_6 = |(in_vaddr >= 64'h80000000 & in_vaddr < 64'h100000000); // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  hasScAccessFault = io__in_valid & _isAmo_T_4 & ~vmEnable & ~_hasScAccessFault_T_6; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 84:58]
  wire  valid = io__in_valid & addrAligned & ~hasScAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 86:39]
  wire  _io_vaddr_T_2 = hasAddrMisaligned | hasScAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 91:44]
  reg [63:0] io_vaddr_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [63:0] _GEN_0 = _io_vaddr_T_2 ? in_vaddr : io_vaddr_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  wire  atomReq = valid & isAtomic; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 97:23]
  wire  amoReq = valid & isAmo; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 98:22]
  wire  lrReq = valid & _isAmo_T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 99:21]
  wire  scReq = valid & _isAmo_T_4; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 100:21]
  wire [2:0] funct3 = io__instr[14:12]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 108:24]
  wire  scInvalid = scReq & (io__in_bits_src1 != lr_addr | ~lr_0) & _hasScAccessFault_T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 126:53]
  reg [2:0] state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 132:22]
  reg [63:0] atomMemReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
  reg [63:0] atomRegReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
  wire  _T = 3'h0 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
  wire  _lsExecUnit_io_in_valid_T = ~atomReq; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 184:48]
  wire  _io_in_ready_T_1 = lsExecUnit_io__out_ready & lsExecUnit_io__out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _GEN_2 = amoReq ? 3'h5 : 3'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 192:15 195:{19,26}]
  wire [2:0] _GEN_3 = lrReq ? 3'h3 : _GEN_2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 196:{18,25}]
  wire [2:0] _state_T = scInvalid ? 3'h0 : 3'h4; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 197:31]
  wire  _T_1 = 3'h1 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
  wire [2:0] _GEN_5 = io__out_valid ? 3'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 132:22 211:{26,33}]
  wire [1:0] _lsExecUnit_io_in_bits_func_T = funct3[0] ? 2'h3 : 2'h2; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 231:40]
  wire [2:0] _GEN_6 = _io_in_ready_T_1 ? 3'h6 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 235:37 236:15 132:22]
  wire [3:0] _lsExecUnit_io_in_bits_func_T_1 = funct3[0] ? 4'hb : 4'ha; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 262:40]
  wire [2:0] _GEN_7 = _io_in_ready_T_1 ? 3'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 266:37 267:15 132:22]
  wire  _io_in_ready_T_7 = ~scIsSuccess_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 292:63]
  wire  _io_in_ready_T_8 = _io_in_ready_T_1 | ~scIsSuccess_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 292:60]
  wire [2:0] _GEN_9 = _io_in_ready_T_8 ? 3'h0 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 294:51 295:15 132:22]
  wire  _GEN_15 = 3'h4 == state & (_io_in_ready_T_1 | ~scIsSuccess_0); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 167:30 292:34]
  wire [2:0] _GEN_17 = 3'h4 == state ? _GEN_9 : state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 132:22]
  wire  _GEN_18 = 3'h3 == state | 3'h4 == state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 272:34]
  wire [3:0] _GEN_21 = 3'h3 == state ? {{2'd0}, _lsExecUnit_io_in_bits_func_T} : _lsExecUnit_io_in_bits_func_T_1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 276:34]
  wire  _GEN_23 = 3'h3 == state ? _io_in_ready_T_1 : _GEN_15; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 278:34]
  wire [2:0] _GEN_25 = 3'h3 == state ? _GEN_7 : _GEN_17; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
  wire  _GEN_26 = 3'h7 == state | _GEN_18; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 258:34]
  wire [3:0] _GEN_29 = 3'h7 == state ? _lsExecUnit_io_in_bits_func_T_1 : _GEN_21; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 262:34]
  wire [63:0] _GEN_30 = 3'h7 == state ? atomMemReg : io__wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 263:34]
  wire  _GEN_31 = 3'h7 == state ? _io_in_ready_T_1 : _GEN_23; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 264:34]
  wire [2:0] _GEN_33 = 3'h7 == state ? _GEN_7 : _GEN_25; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
  wire  _GEN_34 = 3'h6 == state ? 1'h0 : _GEN_26; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 244:34]
  wire  _GEN_35 = 3'h6 == state ? 1'h0 : 1'h1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 245:34]
  wire  _GEN_39 = 3'h6 == state ? 1'h0 : _GEN_31; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 250:34]
  wire [2:0] _GEN_41 = 3'h6 == state ? 3'h7 : _GEN_33; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 252:13]
  wire  _GEN_43 = 3'h5 == state | _GEN_34; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 227:34]
  wire  _GEN_44 = 3'h5 == state | _GEN_35; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 228:34]
  wire [3:0] _GEN_46 = 3'h5 == state ? {{2'd0}, _lsExecUnit_io_in_bits_func_T} : _GEN_29; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 231:34]
  wire  _GEN_48 = 3'h5 == state ? 1'h0 : _GEN_39; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 233:34]
  wire [2:0] _GEN_50 = 3'h5 == state ? _GEN_6 : _GEN_41; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
  wire  _GEN_53 = 3'h1 == state | _GEN_43; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 202:34]
  wire  _GEN_54 = 3'h1 == state | _GEN_44; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 203:34]
  wire [6:0] _GEN_56 = 3'h1 == state ? io__in_bits_func : {{3'd0}, _GEN_46}; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 206:34]
  wire [63:0] _GEN_57 = 3'h1 == state ? io__wdata : _GEN_30; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 207:34]
  wire  _GEN_59 = 3'h1 == state ? lsExecUnit_io__out_valid : _GEN_48; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 209:34]
  wire  _GEN_69 = 3'h0 == state ? lsExecUnit_io__out_valid | scInvalid : _GEN_59; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 191:36]
  wire  _hasException_T_1 = lsExecUnit_io__dtlbAF | lsExecUnit_io__dtlbPF | io__loadAddrMisaligned; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 300:67]
  wire  _hasException_T_3 = _hasException_T_1 | io__storeAddrMisaligned | io__loadAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 301:53]
  wire  hasException = _hasException_T_3 | io__storeAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 302:24]
  wire [31:0] lr_paddr = dtlb_paddr[31:0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 316:26]
  wire  _io_out_bits_T_1 = scInvalid | _io_in_ready_T_7; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 324:39]
  wire [63:0] _io_out_bits_T_3 = state == 3'h7 ? atomRegReg : lsExecUnit_io__out_bits; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 324:59]
  reg  mmioReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 329:24]
  wire  setLr = io__out_valid & (lrReq | scReq); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 318:24]
  wire  setLrVal = lrReq & ~hasException; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 319:21]
  wire [63:0] setLrAddr = vmEnable ? {{32'd0}, lr_paddr} : io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 320:19]
  wire  scInflight = state == 3'h4; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 143:23]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [63:0] io_vaddr_r_p; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [63:0] io_vaddr_r_t = io_vaddr_r ^ io_vaddr_r_p; // @[src/main/scala/utils/Hold.scala 23:65]
  wire  toggle_2936_clock;
  wire  toggle_2936_reset;
  wire [63:0] toggle_2936_valid;
  reg [63:0] toggle_2936_valid_reg;
  reg [2:0] state_p; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 132:22]
  wire [2:0] state_t = state ^ state_p; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 132:22]
  wire  toggle_3000_clock;
  wire  toggle_3000_reset;
  wire [2:0] toggle_3000_valid;
  reg [2:0] toggle_3000_valid_reg;
  reg [63:0] atomMemReg_p; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
  wire [63:0] atomMemReg_t = atomMemReg ^ atomMemReg_p; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
  wire  toggle_3003_clock;
  wire  toggle_3003_reset;
  wire [63:0] toggle_3003_valid;
  reg [63:0] toggle_3003_valid_reg;
  reg [63:0] atomRegReg_p; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
  wire [63:0] atomRegReg_t = atomRegReg ^ atomRegReg_p; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
  wire  toggle_3067_clock;
  wire  toggle_3067_reset;
  wire [63:0] toggle_3067_valid;
  reg [63:0] toggle_3067_valid_reg;
  reg  mmioReg_p; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 329:24]
  wire  mmioReg_t = mmioReg ^ mmioReg_p; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 329:24]
  wire  toggle_3131_clock;
  wire  toggle_3131_reset;
  wire  toggle_3131_valid;
  reg  toggle_3131_valid_reg;
  LSExecUnit lsExecUnit ( // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 88:26]
    .clock(lsExecUnit_clock),
    .reset(lsExecUnit_reset),
    .io__in_ready(lsExecUnit_io__in_ready),
    .io__in_valid(lsExecUnit_io__in_valid),
    .io__in_bits_src1(lsExecUnit_io__in_bits_src1),
    .io__in_bits_func(lsExecUnit_io__in_bits_func),
    .io__out_ready(lsExecUnit_io__out_ready),
    .io__out_valid(lsExecUnit_io__out_valid),
    .io__out_bits(lsExecUnit_io__out_bits),
    .io__wdata(lsExecUnit_io__wdata),
    .io__dmem_req_ready(lsExecUnit_io__dmem_req_ready),
    .io__dmem_req_valid(lsExecUnit_io__dmem_req_valid),
    .io__dmem_req_bits_addr(lsExecUnit_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(lsExecUnit_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(lsExecUnit_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(lsExecUnit_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(lsExecUnit_io__dmem_req_bits_wdata),
    .io__dmem_resp_ready(lsExecUnit_io__dmem_resp_ready),
    .io__dmem_resp_valid(lsExecUnit_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(lsExecUnit_io__dmem_resp_bits_rdata),
    .io__isMMIO(lsExecUnit_io__isMMIO),
    .io__dtlbPF(lsExecUnit_io__dtlbPF),
    .io__dtlbAF(lsExecUnit_io__dtlbAF),
    .io__vaddr(lsExecUnit_io__vaddr),
    .io__loadAccessFault(lsExecUnit_io__loadAccessFault),
    .io__storeAccessFault(lsExecUnit_io__storeAccessFault),
    .DTLBPF(lsExecUnit_DTLBPF),
    .scIsSuccess_0(lsExecUnit_scIsSuccess_0),
    .vmEnable_0(lsExecUnit_vmEnable_0),
    .ISAMO2(lsExecUnit_ISAMO2),
    .DTLBFINISH(lsExecUnit_DTLBFINISH),
    .DTLBAF(lsExecUnit_DTLBAF)
  );
  AtomALU atomALU ( // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 135:23]
    .clock(atomALU_clock),
    .reset(atomALU_reset),
    .io_src1(atomALU_io_src1),
    .io_src2(atomALU_io_src2),
    .io_func(atomALU_io_func),
    .io_isWordOp(atomALU_io_isWordOp),
    .io_result(atomALU_io_result)
  );
  GEN_w64_toggle #(.COVER_INDEX(2936)) toggle_2936 (
    .clock(toggle_2936_clock),
    .reset(toggle_2936_reset),
    .valid(toggle_2936_valid)
  );
  GEN_w3_toggle #(.COVER_INDEX(3000)) toggle_3000 (
    .clock(toggle_3000_clock),
    .reset(toggle_3000_reset),
    .valid(toggle_3000_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(3003)) toggle_3003 (
    .clock(toggle_3003_clock),
    .reset(toggle_3003_reset),
    .valid(toggle_3003_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(3067)) toggle_3067 (
    .clock(toggle_3067_clock),
    .reset(toggle_3067_reset),
    .valid(toggle_3067_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(3131)) toggle_3131 (
    .clock(toggle_3131_clock),
    .reset(toggle_3131_reset),
    .valid(toggle_3131_valid)
  );
  assign io__out_valid = hasException | _GEN_69; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 303:23 305:18]
  assign io__out_bits = scReq ? {{63'd0}, _io_out_bits_T_1} : _io_out_bits_T_3; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 324:21]
  assign io__dmem_req_valid = lsExecUnit_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign io__dmem_req_bits_addr = lsExecUnit_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign io__dmem_req_bits_size = lsExecUnit_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign io__dmem_req_bits_cmd = lsExecUnit_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign io__dmem_req_bits_wmask = lsExecUnit_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign io__dmem_req_bits_wdata = lsExecUnit_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign io__isMMIO = mmioReg & io__out_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 332:24]
  assign io__dtlbPF = lsExecUnit_io__dtlbPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 94:13]
  assign io__dtlbAF = lsExecUnit_io__dtlbAF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 95:13]
  assign io__vaddr = io__loadAddrMisaligned | io__storeAddrMisaligned | hasScAccessFault ? _GEN_0 : lsExecUnit_io__vaddr
    ; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 90:18]
  assign io__loadAddrMisaligned = hasAddrMisaligned & (_io_loadAddrMisaligned_T_4 | _isAmo_T_1); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 74:46]
  assign io__storeAddrMisaligned = hasAddrMisaligned & (io__in_bits_func[3] | isAmo | _isAmo_T_4); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 75:47]
  assign io__loadAccessFault = lsExecUnit_io__loadAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 334:22]
  assign io__storeAccessFault = lsExecUnit_io__storeAccessFault | hasScAccessFault; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 335:57]
  assign setLr_0 = setLr;
  assign scInflight_0 = scInflight;
  assign amoReq_0 = amoReq;
  assign setLrVal_0 = setLrVal;
  assign setLrAddr_0 = setLrAddr;
  assign lsExecUnit_clock = clock;
  assign lsExecUnit_reset = reset;
  assign lsExecUnit_io__in_valid = 3'h0 == state ? valid & ~atomReq : _GEN_53; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 184:36]
  assign lsExecUnit_io__in_bits_src1 = 3'h0 == state ? _in_vaddr_T_1 : io__in_bits_src1; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 186:36]
  assign lsExecUnit_io__in_bits_func = 3'h0 == state ? io__in_bits_func : _GEN_56; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 188:36]
  assign lsExecUnit_io__out_ready = 3'h0 == state | _GEN_54; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 185:36]
  assign lsExecUnit_io__wdata = 3'h0 == state ? io__wdata : _GEN_57; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18 189:36]
  assign lsExecUnit_io__dmem_req_ready = io__dmem_req_ready; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign lsExecUnit_io__dmem_resp_valid = io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign lsExecUnit_io__dmem_resp_bits_rdata = io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 322:11]
  assign lsExecUnit_DTLBPF = _T_12_0;
  assign lsExecUnit_scIsSuccess_0 = scIsSuccess_0;
  assign lsExecUnit_vmEnable_0 = vmEnable;
  assign lsExecUnit_ISAMO2 = amoReq;
  assign lsExecUnit_DTLBFINISH = DTLBFINISH;
  assign lsExecUnit_DTLBAF = _T_13_1;
  assign atomALU_clock = clock;
  assign atomALU_reset = reset;
  assign atomALU_io_src1 = atomMemReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 136:19]
  assign atomALU_io_src2 = io__wdata; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 137:19]
  assign atomALU_io_func = io__in_bits_func; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 138:19]
  assign atomALU_io_isWordOp = ~funct3[0]; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 110:20]
  assign toggle_2936_clock = clock;
  assign toggle_2936_reset = reset;
  assign toggle_2936_valid = io_vaddr_r ^ toggle_2936_valid_reg;
  assign toggle_3000_clock = clock;
  assign toggle_3000_reset = reset;
  assign toggle_3000_valid = state ^ toggle_3000_valid_reg;
  assign toggle_3003_clock = clock;
  assign toggle_3003_reset = reset;
  assign toggle_3003_valid = atomMemReg ^ toggle_3003_valid_reg;
  assign toggle_3067_clock = clock;
  assign toggle_3067_reset = reset;
  assign toggle_3067_valid = atomRegReg ^ toggle_3067_valid_reg;
  assign toggle_3131_clock = clock;
  assign toggle_3131_reset = reset;
  assign toggle_3131_valid = mmioReg ^ toggle_3131_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      io_vaddr_r <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_io_vaddr_T_2) begin // @[src/main/scala/utils/Hold.scala 23:65]
      if (isAtomic) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 62:21]
        io_vaddr_r <= io__in_bits_src1;
      end else begin
        io_vaddr_r <= _in_vaddr_T_1;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 132:22]
      state <= 3'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 132:22]
    end else if (hasException) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 303:23]
      state <= 3'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 304:11]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
      if (scReq) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 197:18]
        state <= _state_T; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 197:25]
      end else begin
        state <= _GEN_3;
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
      state <= _GEN_5;
    end else begin
      state <= _GEN_50;
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
        if (3'h5 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
          atomMemReg <= lsExecUnit_io__out_bits; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 239:18]
        end else if (3'h6 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
          atomMemReg <= atomALU_io_result; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 253:18]
        end
      end
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
        if (3'h5 == state) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 171:18]
          atomRegReg <= lsExecUnit_io__out_bits; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 240:18]
        end
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 329:24]
      mmioReg <= 1'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 329:24]
    end else if (io__out_valid) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 331:23]
      mmioReg <= 1'h0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 331:33]
    end else if (~mmioReg) begin // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 330:19]
      mmioReg <= lsuMMIO_0; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 330:29]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T & _T_1 & ~reset & ~(_lsExecUnit_io_in_valid_T | ~amoReq | ~lrReq | ~scReq)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UnpipelinedLSU.scala:210 assert(!atomReq || !amoReq || !lrReq || !scReq)\n"); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 210:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    io_vaddr_r_p <= io_vaddr_r; // @[src/main/scala/utils/Hold.scala 23:65]
    toggle_2936_valid_reg <= io_vaddr_r;
    state_p <= state; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 132:22]
    toggle_3000_valid_reg <= state;
    atomMemReg_p <= atomMemReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    toggle_3003_valid_reg <= atomMemReg;
    atomRegReg_p <= atomRegReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    toggle_3067_valid_reg <= atomRegReg;
    mmioReg_p <= mmioReg; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 329:24]
    toggle_3131_valid_reg <= mmioReg;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  io_vaddr_r = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[2:0];
  _RAND_2 = {2{`RANDOM}};
  atomMemReg = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  atomRegReg = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  mmioReg = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  io_vaddr_r_p = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  toggle_2936_valid_reg = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  state_p = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  toggle_3000_valid_reg = _RAND_8[2:0];
  _RAND_9 = {2{`RANDOM}};
  atomMemReg_p = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  toggle_3003_valid_reg = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  atomRegReg_p = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  toggle_3067_valid_reg = _RAND_12[63:0];
  _RAND_13 = {1{`RANDOM}};
  mmioReg_p = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  toggle_3131_valid_reg = _RAND_14[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~_T & _T_1 & ~reset) begin
      assert(_lsExecUnit_io_in_valid_T | ~amoReq | ~lrReq | ~scReq); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 210:13]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[0]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[1]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[2]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[3]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[4]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[5]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[6]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[7]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[8]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[9]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[10]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[11]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[12]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[13]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[14]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[15]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[16]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[17]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[18]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[19]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[20]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[21]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[22]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[23]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[24]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[25]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[26]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[27]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[28]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[29]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[30]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[31]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[32]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[33]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[34]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[35]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[36]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[37]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[38]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[39]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[40]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[41]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[42]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[43]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[44]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[45]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[46]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[47]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[48]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[49]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[50]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[51]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[52]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[53]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[54]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[55]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[56]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[57]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[58]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[59]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[60]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[61]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[62]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(io_vaddr_r_t[63]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(state_t[0]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 132:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[1]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 132:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[2]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 132:22]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[0]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[1]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[2]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[3]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[4]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[5]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[6]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[7]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[8]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[9]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[10]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[11]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[12]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[13]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[14]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[15]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[16]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[17]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[18]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[19]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[20]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[21]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[22]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[23]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[24]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[25]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[26]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[27]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[28]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[29]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[30]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[31]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[32]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[33]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[34]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[35]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[36]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[37]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[38]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[39]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[40]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[41]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[42]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[43]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[44]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[45]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[46]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[47]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[48]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[49]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[50]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[51]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[52]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[53]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[54]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[55]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[56]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[57]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[58]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[59]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[60]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[61]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[62]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomMemReg_t[63]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 133:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[0]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[1]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[2]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[3]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[4]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[5]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[6]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[7]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[8]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[9]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[10]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[11]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[12]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[13]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[14]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[15]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[16]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[17]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[18]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[19]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[20]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[21]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[22]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[23]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[24]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[25]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[26]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[27]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[28]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[29]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[30]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[31]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[32]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[33]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[34]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[35]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[36]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[37]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[38]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[39]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[40]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[41]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[42]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[43]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[44]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[45]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[46]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[47]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[48]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[49]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[50]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[51]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[52]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[53]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[54]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[55]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[56]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[57]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[58]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[59]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[60]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[61]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[62]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(atomRegReg_t[63]); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 134:23]
    end
    //
    if (enToggle_past) begin
      cover(mmioReg_t); // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 329:24]
    end
  end
endmodule
module Multiplier(
  input          clock,
  input          reset,
  output         io_in_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  input          io_in_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  input  [64:0]  io_in_bits_0, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  input  [64:0]  io_in_bits_1, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  input          io_out_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  output         io_out_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
  output [129:0] io_out_bits // @[src/main/scala/nutcore/backend/fu/MDU.scala 53:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [159:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [95:0] _RAND_10;
  reg [95:0] _RAND_11;
  reg [95:0] _RAND_12;
  reg [95:0] _RAND_13;
  reg [159:0] _RAND_14;
  reg [159:0] _RAND_15;
  reg [159:0] _RAND_16;
  reg [159:0] _RAND_17;
  reg [159:0] _RAND_18;
  reg [159:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
`endif // RANDOMIZE_REG_INIT
  reg [64:0] mulRes_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  reg [64:0] mulRes_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  reg [129:0] io_out_bits_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
  reg [129:0] io_out_bits_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
  reg [129:0] io_out_bits_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
  reg  io_out_valid_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  reg  io_out_valid_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
  reg  io_out_valid_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
  reg  io_out_valid_REG_3; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
  reg  busy; // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21]
  wire  _GEN_0 = io_in_valid & ~busy | busy; // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21 63:{31,38}]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [64:0] mulRes_REG_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  wire [64:0] mulRes_REG_t = mulRes_REG ^ mulRes_REG_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  wire  toggle_3132_clock;
  wire  toggle_3132_reset;
  wire [64:0] toggle_3132_valid;
  reg [64:0] toggle_3132_valid_reg;
  reg [64:0] mulRes_REG_1_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  wire [64:0] mulRes_REG_1_t = mulRes_REG_1 ^ mulRes_REG_1_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  wire  toggle_3197_clock;
  wire  toggle_3197_reset;
  wire [64:0] toggle_3197_valid;
  reg [64:0] toggle_3197_valid_reg;
  reg [129:0] io_out_bits_REG_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
  wire [129:0] io_out_bits_REG_t = $signed(io_out_bits_REG) ^ $signed(io_out_bits_REG_p); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
  wire  toggle_3262_clock;
  wire  toggle_3262_reset;
  wire [129:0] toggle_3262_valid;
  reg [129:0] toggle_3262_valid_reg;
  reg [129:0] io_out_bits_REG_1_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
  wire [129:0] io_out_bits_REG_1_t = $signed(io_out_bits_REG_1) ^ $signed(io_out_bits_REG_1_p); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
  wire  toggle_3392_clock;
  wire  toggle_3392_reset;
  wire [129:0] toggle_3392_valid;
  reg [129:0] toggle_3392_valid_reg;
  reg [129:0] io_out_bits_REG_2_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
  wire [129:0] io_out_bits_REG_2_t = $signed(io_out_bits_REG_2) ^ $signed(io_out_bits_REG_2_p); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
  wire  toggle_3522_clock;
  wire  toggle_3522_reset;
  wire [129:0] toggle_3522_valid;
  reg [129:0] toggle_3522_valid_reg;
  reg  io_out_valid_REG_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  wire  io_out_valid_REG_t = io_out_valid_REG ^ io_out_valid_REG_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
  wire  toggle_3652_clock;
  wire  toggle_3652_reset;
  wire  toggle_3652_valid;
  reg  toggle_3652_valid_reg;
  reg  io_out_valid_REG_1_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
  wire  io_out_valid_REG_1_t = io_out_valid_REG_1 ^ io_out_valid_REG_1_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
  wire  toggle_3653_clock;
  wire  toggle_3653_reset;
  wire  toggle_3653_valid;
  reg  toggle_3653_valid_reg;
  reg  io_out_valid_REG_2_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
  wire  io_out_valid_REG_2_t = io_out_valid_REG_2 ^ io_out_valid_REG_2_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
  wire  toggle_3654_clock;
  wire  toggle_3654_reset;
  wire  toggle_3654_valid;
  reg  toggle_3654_valid_reg;
  reg  io_out_valid_REG_3_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
  wire  io_out_valid_REG_3_t = io_out_valid_REG_3 ^ io_out_valid_REG_3_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
  wire  toggle_3655_clock;
  wire  toggle_3655_reset;
  wire  toggle_3655_valid;
  reg  toggle_3655_valid_reg;
  reg  busy_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21]
  wire  busy_t = busy ^ busy_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21]
  wire  toggle_3656_clock;
  wire  toggle_3656_reset;
  wire  toggle_3656_valid;
  reg  toggle_3656_valid_reg;
  GEN_w65_toggle #(.COVER_INDEX(3132)) toggle_3132 (
    .clock(toggle_3132_clock),
    .reset(toggle_3132_reset),
    .valid(toggle_3132_valid)
  );
  GEN_w65_toggle #(.COVER_INDEX(3197)) toggle_3197 (
    .clock(toggle_3197_clock),
    .reset(toggle_3197_reset),
    .valid(toggle_3197_valid)
  );
  GEN_w130_toggle #(.COVER_INDEX(3262)) toggle_3262 (
    .clock(toggle_3262_clock),
    .reset(toggle_3262_reset),
    .valid(toggle_3262_valid)
  );
  GEN_w130_toggle #(.COVER_INDEX(3392)) toggle_3392 (
    .clock(toggle_3392_clock),
    .reset(toggle_3392_reset),
    .valid(toggle_3392_valid)
  );
  GEN_w130_toggle #(.COVER_INDEX(3522)) toggle_3522 (
    .clock(toggle_3522_clock),
    .reset(toggle_3522_reset),
    .valid(toggle_3522_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(3652)) toggle_3652 (
    .clock(toggle_3652_clock),
    .reset(toggle_3652_reset),
    .valid(toggle_3652_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(3653)) toggle_3653 (
    .clock(toggle_3653_clock),
    .reset(toggle_3653_reset),
    .valid(toggle_3653_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(3654)) toggle_3654 (
    .clock(toggle_3654_clock),
    .reset(toggle_3654_reset),
    .valid(toggle_3654_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(3655)) toggle_3655 (
    .clock(toggle_3655_clock),
    .reset(toggle_3655_reset),
    .valid(toggle_3655_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(3656)) toggle_3656 (
    .clock(toggle_3656_clock),
    .reset(toggle_3656_reset),
    .valid(toggle_3656_valid)
  );
  assign io_in_ready = ~busy; // @[src/main/scala/nutcore/backend/fu/MDU.scala 65:49]
  assign io_out_valid = io_out_valid_REG_3; // @[src/main/scala/nutcore/backend/fu/MDU.scala 60:16]
  assign io_out_bits = io_out_bits_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 59:37]
  assign toggle_3132_clock = clock;
  assign toggle_3132_reset = reset;
  assign toggle_3132_valid = mulRes_REG ^ toggle_3132_valid_reg;
  assign toggle_3197_clock = clock;
  assign toggle_3197_reset = reset;
  assign toggle_3197_valid = mulRes_REG_1 ^ toggle_3197_valid_reg;
  assign toggle_3262_clock = clock;
  assign toggle_3262_reset = reset;
  assign toggle_3262_valid = $signed(io_out_bits_REG) ^ toggle_3262_valid_reg;
  assign toggle_3392_clock = clock;
  assign toggle_3392_reset = reset;
  assign toggle_3392_valid = $signed(io_out_bits_REG_1) ^ toggle_3392_valid_reg;
  assign toggle_3522_clock = clock;
  assign toggle_3522_reset = reset;
  assign toggle_3522_valid = $signed(io_out_bits_REG_2) ^ toggle_3522_valid_reg;
  assign toggle_3652_clock = clock;
  assign toggle_3652_reset = reset;
  assign toggle_3652_valid = io_out_valid_REG ^ toggle_3652_valid_reg;
  assign toggle_3653_clock = clock;
  assign toggle_3653_reset = reset;
  assign toggle_3653_valid = io_out_valid_REG_1 ^ toggle_3653_valid_reg;
  assign toggle_3654_clock = clock;
  assign toggle_3654_reset = reset;
  assign toggle_3654_valid = io_out_valid_REG_2 ^ toggle_3654_valid_reg;
  assign toggle_3655_clock = clock;
  assign toggle_3655_reset = reset;
  assign toggle_3655_valid = io_out_valid_REG_3 ^ toggle_3655_valid_reg;
  assign toggle_3656_clock = clock;
  assign toggle_3656_reset = reset;
  assign toggle_3656_valid = busy ^ toggle_3656_valid_reg;
  always @(posedge clock) begin
    mulRes_REG <= io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    mulRes_REG_1 <= io_in_bits_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    io_out_bits_REG <= $signed(mulRes_REG) * $signed(mulRes_REG_1); // @[src/main/scala/nutcore/backend/fu/MDU.scala 58:49]
    io_out_bits_REG_1 <= io_out_bits_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    io_out_bits_REG_2 <= io_out_bits_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    io_out_valid_REG <= io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
    io_out_valid_REG_1 <= io_out_valid_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    io_out_valid_REG_2 <= io_out_valid_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    io_out_valid_REG_3 <= io_out_valid_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21]
      busy <= 1'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21]
    end else if (io_out_valid) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 64:23]
      busy <= 1'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 64:30]
    end else begin
      busy <= _GEN_0;
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    mulRes_REG_p <= mulRes_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    toggle_3132_valid_reg <= mulRes_REG;
    mulRes_REG_1_p <= mulRes_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    toggle_3197_valid_reg <= mulRes_REG_1;
    io_out_bits_REG_p <= io_out_bits_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    toggle_3262_valid_reg <= io_out_bits_REG;
    io_out_bits_REG_1_p <= io_out_bits_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    toggle_3392_valid_reg <= io_out_bits_REG_1;
    io_out_bits_REG_2_p <= io_out_bits_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    toggle_3522_valid_reg <= io_out_bits_REG_2;
    io_out_valid_REG_p <= io_out_valid_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    toggle_3652_valid_reg <= io_out_valid_REG;
    io_out_valid_REG_1_p <= io_out_valid_REG_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    toggle_3653_valid_reg <= io_out_valid_REG_1;
    io_out_valid_REG_2_p <= io_out_valid_REG_2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    toggle_3654_valid_reg <= io_out_valid_REG_2;
    io_out_valid_REG_3_p <= io_out_valid_REG_3; // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    toggle_3655_valid_reg <= io_out_valid_REG_3;
    busy_p <= busy; // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21]
    toggle_3656_valid_reg <= busy;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  mulRes_REG = _RAND_0[64:0];
  _RAND_1 = {3{`RANDOM}};
  mulRes_REG_1 = _RAND_1[64:0];
  _RAND_2 = {5{`RANDOM}};
  io_out_bits_REG = _RAND_2[129:0];
  _RAND_3 = {5{`RANDOM}};
  io_out_bits_REG_1 = _RAND_3[129:0];
  _RAND_4 = {5{`RANDOM}};
  io_out_bits_REG_2 = _RAND_4[129:0];
  _RAND_5 = {1{`RANDOM}};
  io_out_valid_REG = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  io_out_valid_REG_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  io_out_valid_REG_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  io_out_valid_REG_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  busy = _RAND_9[0:0];
  _RAND_10 = {3{`RANDOM}};
  mulRes_REG_p = _RAND_10[64:0];
  _RAND_11 = {3{`RANDOM}};
  toggle_3132_valid_reg = _RAND_11[64:0];
  _RAND_12 = {3{`RANDOM}};
  mulRes_REG_1_p = _RAND_12[64:0];
  _RAND_13 = {3{`RANDOM}};
  toggle_3197_valid_reg = _RAND_13[64:0];
  _RAND_14 = {5{`RANDOM}};
  io_out_bits_REG_p = _RAND_14[129:0];
  _RAND_15 = {5{`RANDOM}};
  toggle_3262_valid_reg = _RAND_15[129:0];
  _RAND_16 = {5{`RANDOM}};
  io_out_bits_REG_1_p = _RAND_16[129:0];
  _RAND_17 = {5{`RANDOM}};
  toggle_3392_valid_reg = _RAND_17[129:0];
  _RAND_18 = {5{`RANDOM}};
  io_out_bits_REG_2_p = _RAND_18[129:0];
  _RAND_19 = {5{`RANDOM}};
  toggle_3522_valid_reg = _RAND_19[129:0];
  _RAND_20 = {1{`RANDOM}};
  io_out_valid_REG_p = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  toggle_3652_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  io_out_valid_REG_1_p = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  toggle_3653_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  io_out_valid_REG_2_p = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  toggle_3654_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  io_out_valid_REG_3_p = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  toggle_3655_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  busy_p = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  toggle_3656_valid_reg = _RAND_29[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[0]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[1]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[2]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[3]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[4]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[5]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[6]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[7]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[8]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[9]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[10]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[11]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[12]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[13]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[14]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[15]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[16]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[17]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[18]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[19]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[20]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[21]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[22]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[23]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[24]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[25]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[26]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[27]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[28]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[29]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[30]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[31]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[32]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[33]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[34]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[35]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[36]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[37]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[38]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[39]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[40]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[41]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[42]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[43]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[44]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[45]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[46]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[47]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[48]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[49]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[50]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[51]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[52]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[53]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[54]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[55]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[56]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[57]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[58]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[59]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[60]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[61]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[62]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[63]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_t[64]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[0]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[1]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[2]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[3]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[4]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[5]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[6]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[7]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[8]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[9]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[10]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[11]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[12]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[13]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[14]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[15]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[16]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[17]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[18]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[19]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[20]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[21]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[22]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[23]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[24]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[25]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[26]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[27]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[28]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[29]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[30]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[31]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[32]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[33]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[34]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[35]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[36]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[37]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[38]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[39]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[40]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[41]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[42]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[43]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[44]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[45]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[46]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[47]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[48]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[49]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[50]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[51]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[52]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[53]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[54]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[55]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[56]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[57]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[58]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[59]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[60]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[61]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[62]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[63]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(mulRes_REG_1_t[64]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[0]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[1]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[2]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[3]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[4]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[5]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[6]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[7]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[8]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[9]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[10]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[11]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[12]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[13]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[14]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[15]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[16]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[17]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[18]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[19]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[20]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[21]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[22]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[23]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[24]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[25]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[26]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[27]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[28]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[29]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[30]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[31]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[32]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[33]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[34]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[35]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[36]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[37]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[38]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[39]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[40]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[41]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[42]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[43]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[44]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[45]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[46]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[47]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[48]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[49]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[50]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[51]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[52]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[53]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[54]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[55]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[56]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[57]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[58]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[59]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[60]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[61]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[62]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[63]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[64]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[65]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[66]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[67]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[68]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[69]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[70]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[71]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[72]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[73]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[74]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[75]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[76]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[77]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[78]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[79]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[80]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[81]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[82]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[83]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[84]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[85]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[86]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[87]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[88]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[89]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[90]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[91]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[92]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[93]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[94]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[95]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[96]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[97]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[98]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[99]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[100]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[101]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[102]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[103]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[104]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[105]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[106]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[107]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[108]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[109]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[110]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[111]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[112]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[113]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[114]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[115]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[116]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[117]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[118]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[119]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[120]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[121]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[122]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[123]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[124]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[125]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[126]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[127]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[128]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_t[129]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[0]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[1]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[2]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[3]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[4]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[5]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[6]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[7]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[8]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[9]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[10]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[11]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[12]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[13]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[14]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[15]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[16]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[17]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[18]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[19]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[20]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[21]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[22]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[23]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[24]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[25]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[26]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[27]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[28]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[29]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[30]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[31]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[32]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[33]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[34]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[35]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[36]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[37]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[38]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[39]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[40]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[41]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[42]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[43]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[44]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[45]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[46]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[47]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[48]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[49]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[50]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[51]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[52]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[53]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[54]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[55]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[56]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[57]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[58]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[59]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[60]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[61]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[62]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[63]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[64]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[65]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[66]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[67]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[68]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[69]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[70]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[71]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[72]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[73]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[74]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[75]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[76]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[77]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[78]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[79]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[80]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[81]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[82]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[83]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[84]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[85]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[86]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[87]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[88]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[89]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[90]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[91]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[92]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[93]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[94]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[95]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[96]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[97]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[98]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[99]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[100]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[101]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[102]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[103]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[104]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[105]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[106]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[107]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[108]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[109]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[110]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[111]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[112]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[113]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[114]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[115]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[116]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[117]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[118]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[119]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[120]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[121]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[122]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[123]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[124]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[125]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[126]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[127]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[128]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_1_t[129]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[0]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[1]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[2]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[3]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[4]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[5]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[6]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[7]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[8]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[9]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[10]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[11]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[12]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[13]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[14]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[15]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[16]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[17]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[18]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[19]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[20]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[21]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[22]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[23]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[24]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[25]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[26]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[27]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[28]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[29]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[30]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[31]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[32]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[33]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[34]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[35]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[36]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[37]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[38]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[39]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[40]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[41]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[42]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[43]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[44]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[45]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[46]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[47]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[48]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[49]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[50]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[51]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[52]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[53]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[54]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[55]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[56]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[57]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[58]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[59]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[60]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[61]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[62]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[63]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[64]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[65]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[66]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[67]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[68]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[69]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[70]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[71]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[72]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[73]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[74]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[75]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[76]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[77]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[78]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[79]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[80]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[81]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[82]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[83]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[84]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[85]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[86]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[87]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[88]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[89]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[90]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[91]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[92]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[93]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[94]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[95]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[96]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[97]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[98]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[99]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[100]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[101]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[102]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[103]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[104]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[105]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[106]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[107]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[108]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[109]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[110]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[111]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[112]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[113]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[114]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[115]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[116]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[117]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[118]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[119]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[120]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[121]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[122]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[123]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[124]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[125]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[126]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[127]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[128]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_bits_REG_2_t[129]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(io_out_valid_REG_t); // @[src/main/scala/nutcore/backend/fu/MDU.scala 56:43]
    end
    //
    if (enToggle_past) begin
      cover(io_out_valid_REG_1_t); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:60]
    end
    //
    if (enToggle_past) begin
      cover(io_out_valid_REG_2_t); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:52]
    end
    //
    if (enToggle_past) begin
      cover(io_out_valid_REG_3_t); // @[src/main/scala/nutcore/backend/fu/MDU.scala 57:44]
    end
    //
    if (enToggle_past) begin
      cover(busy_t); // @[src/main/scala/nutcore/backend/fu/MDU.scala 62:21]
    end
  end
endmodule
module Divider(
  input          clock,
  input          reset,
  output         io_in_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  input          io_in_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  input  [63:0]  io_in_bits_0, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  input  [63:0]  io_in_bits_1, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  input          io_sign, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  output         io_out_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
  output [127:0] io_out_bits // @[src/main/scala/nutcore/backend/fu/MDU.scala 69:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [159:0] _RAND_9;
  reg [159:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [95:0] _RAND_17;
  reg [95:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
  wire  _newReq_T_1 = io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  newReq = state == 3'h0 & _newReq_T_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 78:35]
  wire  divBy0 = io_in_bits_1 == 64'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 81:18]
  reg [128:0] shiftReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
  wire [64:0] hi = shiftReg[128:64]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 84:20]
  wire [63:0] lo = shiftReg[63:0]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 85:20]
  wire  aSign = io_in_bits_0[63] & io_sign; // @[src/main/scala/nutcore/backend/fu/MDU.scala 72:24]
  wire [63:0] _T_1 = 64'h0 - io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 73:16]
  wire [63:0] aVal = aSign ? _T_1 : io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 73:12]
  wire  bSign = io_in_bits_1[63] & io_sign; // @[src/main/scala/nutcore/backend/fu/MDU.scala 72:24]
  wire [63:0] _T_3 = 64'h0 - io_in_bits_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 73:16]
  reg  aSignReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 89:27]
  reg  qSignReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 90:27]
  reg [63:0] bReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
  wire [64:0] _aValx2Reg_T = {aVal,1'h0}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:32]
  reg [64:0] aValx2Reg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
  reg [5:0] cnt_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [31:0] canSkipShift_hi = bReg[63:32]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [31:0] canSkipShift_lo = bReg[31:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi = |canSkipShift_hi; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [15:0] canSkipShift_hi_1 = canSkipShift_hi[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] canSkipShift_lo_1 = canSkipShift_hi[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_1 = |canSkipShift_hi_1; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] canSkipShift_hi_2 = canSkipShift_hi_1[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_2 = canSkipShift_hi_1[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_2 = |canSkipShift_hi_2; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_3 = canSkipShift_hi_2[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_3 = canSkipShift_hi_2[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_3 = |canSkipShift_hi_3; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_3 = canSkipShift_hi_3[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_3[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_4 = canSkipShift_hi_3[3] ? 2'h3 : _canSkipShift_T_3; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_8 = canSkipShift_lo_3[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_3[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_9 = canSkipShift_lo_3[3] ? 2'h3 : _canSkipShift_T_8; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_10 = canSkipShift_useHi_3 ? _canSkipShift_T_4 : _canSkipShift_T_9; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_11 = {canSkipShift_useHi_3,_canSkipShift_T_10}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_4 = canSkipShift_lo_2[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_4 = canSkipShift_lo_2[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_4 = |canSkipShift_hi_4; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_15 = canSkipShift_hi_4[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_4[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_16 = canSkipShift_hi_4[3] ? 2'h3 : _canSkipShift_T_15; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_20 = canSkipShift_lo_4[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_4[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_21 = canSkipShift_lo_4[3] ? 2'h3 : _canSkipShift_T_20; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_22 = canSkipShift_useHi_4 ? _canSkipShift_T_16 : _canSkipShift_T_21; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_23 = {canSkipShift_useHi_4,_canSkipShift_T_22}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_24 = canSkipShift_useHi_2 ? _canSkipShift_T_11 : _canSkipShift_T_23; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_25 = {canSkipShift_useHi_2,_canSkipShift_T_24}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] canSkipShift_hi_5 = canSkipShift_lo_1[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_5 = canSkipShift_lo_1[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_5 = |canSkipShift_hi_5; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_6 = canSkipShift_hi_5[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_6 = canSkipShift_hi_5[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_6 = |canSkipShift_hi_6; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_29 = canSkipShift_hi_6[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_6[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_30 = canSkipShift_hi_6[3] ? 2'h3 : _canSkipShift_T_29; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_34 = canSkipShift_lo_6[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_6[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_35 = canSkipShift_lo_6[3] ? 2'h3 : _canSkipShift_T_34; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_36 = canSkipShift_useHi_6 ? _canSkipShift_T_30 : _canSkipShift_T_35; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_37 = {canSkipShift_useHi_6,_canSkipShift_T_36}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_7 = canSkipShift_lo_5[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_7 = canSkipShift_lo_5[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_7 = |canSkipShift_hi_7; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_41 = canSkipShift_hi_7[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_7[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_42 = canSkipShift_hi_7[3] ? 2'h3 : _canSkipShift_T_41; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_46 = canSkipShift_lo_7[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_7[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_47 = canSkipShift_lo_7[3] ? 2'h3 : _canSkipShift_T_46; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_48 = canSkipShift_useHi_7 ? _canSkipShift_T_42 : _canSkipShift_T_47; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_49 = {canSkipShift_useHi_7,_canSkipShift_T_48}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_50 = canSkipShift_useHi_5 ? _canSkipShift_T_37 : _canSkipShift_T_49; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_51 = {canSkipShift_useHi_5,_canSkipShift_T_50}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _canSkipShift_T_52 = canSkipShift_useHi_1 ? _canSkipShift_T_25 : _canSkipShift_T_51; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _canSkipShift_T_53 = {canSkipShift_useHi_1,_canSkipShift_T_52}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [15:0] canSkipShift_hi_8 = canSkipShift_lo[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] canSkipShift_lo_8 = canSkipShift_lo[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_8 = |canSkipShift_hi_8; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] canSkipShift_hi_9 = canSkipShift_hi_8[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_9 = canSkipShift_hi_8[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_9 = |canSkipShift_hi_9; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_10 = canSkipShift_hi_9[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_10 = canSkipShift_hi_9[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_10 = |canSkipShift_hi_10; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_57 = canSkipShift_hi_10[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_10[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_58 = canSkipShift_hi_10[3] ? 2'h3 : _canSkipShift_T_57; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_62 = canSkipShift_lo_10[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_10[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_63 = canSkipShift_lo_10[3] ? 2'h3 : _canSkipShift_T_62; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_64 = canSkipShift_useHi_10 ? _canSkipShift_T_58 : _canSkipShift_T_63; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_65 = {canSkipShift_useHi_10,_canSkipShift_T_64}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_11 = canSkipShift_lo_9[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_11 = canSkipShift_lo_9[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_11 = |canSkipShift_hi_11; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_69 = canSkipShift_hi_11[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_11[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_70 = canSkipShift_hi_11[3] ? 2'h3 : _canSkipShift_T_69; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_74 = canSkipShift_lo_11[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_11[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_75 = canSkipShift_lo_11[3] ? 2'h3 : _canSkipShift_T_74; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_76 = canSkipShift_useHi_11 ? _canSkipShift_T_70 : _canSkipShift_T_75; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_77 = {canSkipShift_useHi_11,_canSkipShift_T_76}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_78 = canSkipShift_useHi_9 ? _canSkipShift_T_65 : _canSkipShift_T_77; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_79 = {canSkipShift_useHi_9,_canSkipShift_T_78}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] canSkipShift_hi_12 = canSkipShift_lo_8[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_12 = canSkipShift_lo_8[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_12 = |canSkipShift_hi_12; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_13 = canSkipShift_hi_12[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_13 = canSkipShift_hi_12[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_13 = |canSkipShift_hi_13; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_83 = canSkipShift_hi_13[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_13[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_84 = canSkipShift_hi_13[3] ? 2'h3 : _canSkipShift_T_83; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_88 = canSkipShift_lo_13[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_13[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_89 = canSkipShift_lo_13[3] ? 2'h3 : _canSkipShift_T_88; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_90 = canSkipShift_useHi_13 ? _canSkipShift_T_84 : _canSkipShift_T_89; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_91 = {canSkipShift_useHi_13,_canSkipShift_T_90}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_14 = canSkipShift_lo_12[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_14 = canSkipShift_lo_12[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_14 = |canSkipShift_hi_14; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_95 = canSkipShift_hi_14[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_14[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_96 = canSkipShift_hi_14[3] ? 2'h3 : _canSkipShift_T_95; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_100 = canSkipShift_lo_14[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_14[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_101 = canSkipShift_lo_14[3] ? 2'h3 : _canSkipShift_T_100; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_102 = canSkipShift_useHi_14 ? _canSkipShift_T_96 : _canSkipShift_T_101; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_103 = {canSkipShift_useHi_14,_canSkipShift_T_102}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_104 = canSkipShift_useHi_12 ? _canSkipShift_T_91 : _canSkipShift_T_103; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_105 = {canSkipShift_useHi_12,_canSkipShift_T_104}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _canSkipShift_T_106 = canSkipShift_useHi_8 ? _canSkipShift_T_79 : _canSkipShift_T_105; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _canSkipShift_T_107 = {canSkipShift_useHi_8,_canSkipShift_T_106}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [4:0] _canSkipShift_T_108 = canSkipShift_useHi ? _canSkipShift_T_53 : _canSkipShift_T_107; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [5:0] _canSkipShift_T_109 = {canSkipShift_useHi,_canSkipShift_T_108}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [6:0] _GEN_20 = {{1'd0}, _canSkipShift_T_109}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 105:31]
  wire [6:0] _canSkipShift_T_110 = 7'h40 | _GEN_20; // @[src/main/scala/nutcore/backend/fu/MDU.scala 105:31]
  wire  canSkipShift_hi_15 = aValx2Reg[64]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [63:0] canSkipShift_lo_15 = aValx2Reg[63:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_15 = |canSkipShift_hi_15; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [31:0] canSkipShift_hi_16 = canSkipShift_lo_15[63:32]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [31:0] canSkipShift_lo_16 = canSkipShift_lo_15[31:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_16 = |canSkipShift_hi_16; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [15:0] canSkipShift_hi_17 = canSkipShift_hi_16[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] canSkipShift_lo_17 = canSkipShift_hi_16[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_17 = |canSkipShift_hi_17; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] canSkipShift_hi_18 = canSkipShift_hi_17[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_18 = canSkipShift_hi_17[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_18 = |canSkipShift_hi_18; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_19 = canSkipShift_hi_18[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_19 = canSkipShift_hi_18[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_19 = |canSkipShift_hi_19; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_114 = canSkipShift_hi_19[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_19[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_115 = canSkipShift_hi_19[3] ? 2'h3 : _canSkipShift_T_114; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_119 = canSkipShift_lo_19[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_19[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_120 = canSkipShift_lo_19[3] ? 2'h3 : _canSkipShift_T_119; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_121 = canSkipShift_useHi_19 ? _canSkipShift_T_115 : _canSkipShift_T_120; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_122 = {canSkipShift_useHi_19,_canSkipShift_T_121}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_20 = canSkipShift_lo_18[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_20 = canSkipShift_lo_18[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_20 = |canSkipShift_hi_20; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_126 = canSkipShift_hi_20[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_20[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_127 = canSkipShift_hi_20[3] ? 2'h3 : _canSkipShift_T_126; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_131 = canSkipShift_lo_20[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_20[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_132 = canSkipShift_lo_20[3] ? 2'h3 : _canSkipShift_T_131; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_133 = canSkipShift_useHi_20 ? _canSkipShift_T_127 : _canSkipShift_T_132; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_134 = {canSkipShift_useHi_20,_canSkipShift_T_133}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_135 = canSkipShift_useHi_18 ? _canSkipShift_T_122 : _canSkipShift_T_134; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_136 = {canSkipShift_useHi_18,_canSkipShift_T_135}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] canSkipShift_hi_21 = canSkipShift_lo_17[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_21 = canSkipShift_lo_17[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_21 = |canSkipShift_hi_21; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_22 = canSkipShift_hi_21[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_22 = canSkipShift_hi_21[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_22 = |canSkipShift_hi_22; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_140 = canSkipShift_hi_22[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_22[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_141 = canSkipShift_hi_22[3] ? 2'h3 : _canSkipShift_T_140; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_145 = canSkipShift_lo_22[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_22[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_146 = canSkipShift_lo_22[3] ? 2'h3 : _canSkipShift_T_145; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_147 = canSkipShift_useHi_22 ? _canSkipShift_T_141 : _canSkipShift_T_146; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_148 = {canSkipShift_useHi_22,_canSkipShift_T_147}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_23 = canSkipShift_lo_21[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_23 = canSkipShift_lo_21[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_23 = |canSkipShift_hi_23; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_152 = canSkipShift_hi_23[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_23[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_153 = canSkipShift_hi_23[3] ? 2'h3 : _canSkipShift_T_152; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_157 = canSkipShift_lo_23[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_23[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_158 = canSkipShift_lo_23[3] ? 2'h3 : _canSkipShift_T_157; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_159 = canSkipShift_useHi_23 ? _canSkipShift_T_153 : _canSkipShift_T_158; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_160 = {canSkipShift_useHi_23,_canSkipShift_T_159}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_161 = canSkipShift_useHi_21 ? _canSkipShift_T_148 : _canSkipShift_T_160; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_162 = {canSkipShift_useHi_21,_canSkipShift_T_161}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _canSkipShift_T_163 = canSkipShift_useHi_17 ? _canSkipShift_T_136 : _canSkipShift_T_162; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _canSkipShift_T_164 = {canSkipShift_useHi_17,_canSkipShift_T_163}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [15:0] canSkipShift_hi_24 = canSkipShift_lo_16[31:16]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [15:0] canSkipShift_lo_24 = canSkipShift_lo_16[15:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_24 = |canSkipShift_hi_24; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [7:0] canSkipShift_hi_25 = canSkipShift_hi_24[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_25 = canSkipShift_hi_24[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_25 = |canSkipShift_hi_25; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_26 = canSkipShift_hi_25[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_26 = canSkipShift_hi_25[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_26 = |canSkipShift_hi_26; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_168 = canSkipShift_hi_26[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_26[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_169 = canSkipShift_hi_26[3] ? 2'h3 : _canSkipShift_T_168; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_173 = canSkipShift_lo_26[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_26[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_174 = canSkipShift_lo_26[3] ? 2'h3 : _canSkipShift_T_173; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_175 = canSkipShift_useHi_26 ? _canSkipShift_T_169 : _canSkipShift_T_174; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_176 = {canSkipShift_useHi_26,_canSkipShift_T_175}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_27 = canSkipShift_lo_25[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_27 = canSkipShift_lo_25[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_27 = |canSkipShift_hi_27; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_180 = canSkipShift_hi_27[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_27[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_181 = canSkipShift_hi_27[3] ? 2'h3 : _canSkipShift_T_180; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_185 = canSkipShift_lo_27[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_27[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_186 = canSkipShift_lo_27[3] ? 2'h3 : _canSkipShift_T_185; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_187 = canSkipShift_useHi_27 ? _canSkipShift_T_181 : _canSkipShift_T_186; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_188 = {canSkipShift_useHi_27,_canSkipShift_T_187}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_189 = canSkipShift_useHi_25 ? _canSkipShift_T_176 : _canSkipShift_T_188; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_190 = {canSkipShift_useHi_25,_canSkipShift_T_189}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [7:0] canSkipShift_hi_28 = canSkipShift_lo_24[15:8]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [7:0] canSkipShift_lo_28 = canSkipShift_lo_24[7:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_28 = |canSkipShift_hi_28; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [3:0] canSkipShift_hi_29 = canSkipShift_hi_28[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_29 = canSkipShift_hi_28[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_29 = |canSkipShift_hi_29; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_194 = canSkipShift_hi_29[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_29[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_195 = canSkipShift_hi_29[3] ? 2'h3 : _canSkipShift_T_194; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_199 = canSkipShift_lo_29[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_29[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_200 = canSkipShift_lo_29[3] ? 2'h3 : _canSkipShift_T_199; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_201 = canSkipShift_useHi_29 ? _canSkipShift_T_195 : _canSkipShift_T_200; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_202 = {canSkipShift_useHi_29,_canSkipShift_T_201}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] canSkipShift_hi_30 = canSkipShift_lo_28[7:4]; // @[src/main/scala/chisel3/util/CircuitMath.scala 33:17]
  wire [3:0] canSkipShift_lo_30 = canSkipShift_lo_28[3:0]; // @[src/main/scala/chisel3/util/CircuitMath.scala 34:17]
  wire  canSkipShift_useHi_30 = |canSkipShift_hi_30; // @[src/main/scala/chisel3/util/CircuitMath.scala 35:22]
  wire [1:0] _canSkipShift_T_206 = canSkipShift_hi_30[2] ? 2'h2 : {{1'd0}, canSkipShift_hi_30[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_207 = canSkipShift_hi_30[3] ? 2'h3 : _canSkipShift_T_206; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_211 = canSkipShift_lo_30[2] ? 2'h2 : {{1'd0}, canSkipShift_lo_30[1]}; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_212 = canSkipShift_lo_30[3] ? 2'h3 : _canSkipShift_T_211; // @[src/main/scala/chisel3/util/CircuitMath.scala 30:10]
  wire [1:0] _canSkipShift_T_213 = canSkipShift_useHi_30 ? _canSkipShift_T_207 : _canSkipShift_T_212; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [2:0] _canSkipShift_T_214 = {canSkipShift_useHi_30,_canSkipShift_T_213}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [2:0] _canSkipShift_T_215 = canSkipShift_useHi_28 ? _canSkipShift_T_202 : _canSkipShift_T_214; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [3:0] _canSkipShift_T_216 = {canSkipShift_useHi_28,_canSkipShift_T_215}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [3:0] _canSkipShift_T_217 = canSkipShift_useHi_24 ? _canSkipShift_T_190 : _canSkipShift_T_216; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [4:0] _canSkipShift_T_218 = {canSkipShift_useHi_24,_canSkipShift_T_217}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [4:0] _canSkipShift_T_219 = canSkipShift_useHi_16 ? _canSkipShift_T_164 : _canSkipShift_T_218; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [5:0] _canSkipShift_T_220 = {canSkipShift_useHi_16,_canSkipShift_T_219}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [5:0] _canSkipShift_T_221 = canSkipShift_useHi_15 ? 6'h0 : _canSkipShift_T_220; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:21]
  wire [6:0] _canSkipShift_T_222 = {canSkipShift_useHi_15,_canSkipShift_T_221}; // @[src/main/scala/chisel3/util/CircuitMath.scala 36:10]
  wire [6:0] canSkipShift = _canSkipShift_T_110 - _canSkipShift_T_222; // @[src/main/scala/nutcore/backend/fu/MDU.scala 105:45]
  wire [6:0] _value_T_1 = canSkipShift >= 7'h3f ? 7'h3f : canSkipShift; // @[src/main/scala/nutcore/backend/fu/MDU.scala 109:38]
  wire [6:0] _value_T_2 = divBy0 ? 7'h0 : _value_T_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 109:21]
  wire [127:0] _GEN_24 = {{63'd0}, aValx2Reg}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 112:27]
  wire [127:0] _shiftReg_T = _GEN_24 << cnt_value; // @[src/main/scala/nutcore/backend/fu/MDU.scala 112:27]
  wire [64:0] _GEN_21 = {{1'd0}, bReg}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 115:28]
  wire  enough = hi >= _GEN_21; // @[src/main/scala/nutcore/backend/fu/MDU.scala 115:28]
  wire [64:0] _GEN_22 = {{1'd0}, bReg}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:36]
  wire [64:0] _shiftReg_T_2 = hi - _GEN_22; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:36]
  wire [64:0] _shiftReg_T_3 = enough ? _shiftReg_T_2 : hi; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:24]
  wire [128:0] _shiftReg_T_5 = {_shiftReg_T_3[63:0],lo,enough}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:20]
  wire  wrap = cnt_value == 6'h3f; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [5:0] _value_T_4 = cnt_value + 6'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [2:0] _GEN_4 = wrap ? 3'h4 : state; // @[src/main/scala/nutcore/backend/fu/MDU.scala 118:{36,44} 77:22]
  wire [2:0] _GEN_5 = state == 3'h4 ? 3'h0 : state; // @[src/main/scala/nutcore/backend/fu/MDU.scala 119:36 120:11 77:22]
  wire [5:0] _GEN_7 = state == 3'h3 ? _value_T_4 : cnt_value; // @[src/main/scala/nutcore/backend/fu/MDU.scala 114:37 src/main/scala/chisel3/util/Counter.scala 77:15 61:40]
  wire [2:0] _GEN_8 = state == 3'h3 ? _GEN_4 : _GEN_5; // @[src/main/scala/nutcore/backend/fu/MDU.scala 114:37]
  wire [5:0] _GEN_11 = state == 3'h2 ? cnt_value : _GEN_7; // @[src/main/scala/nutcore/backend/fu/MDU.scala 111:35 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [6:0] _GEN_12 = state == 3'h1 ? _value_T_2 : {{1'd0}, _GEN_11}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 109:15 97:34]
  wire [6:0] _GEN_16 = newReq ? {{1'd0}, cnt_value} : _GEN_12; // @[src/main/scala/nutcore/backend/fu/MDU.scala 95:17 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [63:0] r = hi[64:1]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 123:13]
  wire [63:0] _resQ_T_1 = 64'h0 - lo; // @[src/main/scala/nutcore/backend/fu/MDU.scala 124:28]
  wire [63:0] resQ = qSignReg ? _resQ_T_1 : lo; // @[src/main/scala/nutcore/backend/fu/MDU.scala 124:17]
  wire [63:0] _resR_T_1 = 64'h0 - r; // @[src/main/scala/nutcore/backend/fu/MDU.scala 125:28]
  wire [63:0] resR = aSignReg ? _resR_T_1 : r; // @[src/main/scala/nutcore/backend/fu/MDU.scala 125:17]
  wire [6:0] _GEN_23 = reset ? 7'h0 : _GEN_16; // @[src/main/scala/chisel3/util/Counter.scala 61:{40,40}]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [2:0] state_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
  wire [2:0] state_t = state ^ state_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
  wire  toggle_3657_clock;
  wire  toggle_3657_reset;
  wire [2:0] toggle_3657_valid;
  reg [2:0] toggle_3657_valid_reg;
  reg [128:0] shiftReg_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
  wire [128:0] shiftReg_t = shiftReg ^ shiftReg_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
  wire  toggle_3660_clock;
  wire  toggle_3660_reset;
  wire [128:0] toggle_3660_valid;
  reg [128:0] toggle_3660_valid_reg;
  reg  aSignReg_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 89:27]
  wire  aSignReg_t = aSignReg ^ aSignReg_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 89:27]
  wire  toggle_3789_clock;
  wire  toggle_3789_reset;
  wire  toggle_3789_valid;
  reg  toggle_3789_valid_reg;
  reg  qSignReg_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 90:27]
  wire  qSignReg_t = qSignReg ^ qSignReg_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 90:27]
  wire  toggle_3790_clock;
  wire  toggle_3790_reset;
  wire  toggle_3790_valid;
  reg  toggle_3790_valid_reg;
  reg [63:0] bReg_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
  wire [63:0] bReg_t = bReg ^ bReg_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
  wire  toggle_3791_clock;
  wire  toggle_3791_reset;
  wire [63:0] toggle_3791_valid;
  reg [63:0] toggle_3791_valid_reg;
  reg [64:0] aValx2Reg_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
  wire [64:0] aValx2Reg_t = aValx2Reg ^ aValx2Reg_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
  wire  toggle_3855_clock;
  wire  toggle_3855_reset;
  wire [64:0] toggle_3855_valid;
  reg [64:0] toggle_3855_valid_reg;
  reg [5:0] cnt_value_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [5:0] cnt_value_t = cnt_value ^ cnt_value_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  toggle_3920_clock;
  wire  toggle_3920_reset;
  wire [5:0] toggle_3920_valid;
  reg [5:0] toggle_3920_valid_reg;
  GEN_w3_toggle #(.COVER_INDEX(3657)) toggle_3657 (
    .clock(toggle_3657_clock),
    .reset(toggle_3657_reset),
    .valid(toggle_3657_valid)
  );
  GEN_w129_toggle #(.COVER_INDEX(3660)) toggle_3660 (
    .clock(toggle_3660_clock),
    .reset(toggle_3660_reset),
    .valid(toggle_3660_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(3789)) toggle_3789 (
    .clock(toggle_3789_clock),
    .reset(toggle_3789_reset),
    .valid(toggle_3789_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(3790)) toggle_3790 (
    .clock(toggle_3790_clock),
    .reset(toggle_3790_reset),
    .valid(toggle_3790_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(3791)) toggle_3791 (
    .clock(toggle_3791_clock),
    .reset(toggle_3791_reset),
    .valid(toggle_3791_valid)
  );
  GEN_w65_toggle #(.COVER_INDEX(3855)) toggle_3855 (
    .clock(toggle_3855_clock),
    .reset(toggle_3855_reset),
    .valid(toggle_3855_valid)
  );
  GEN_w6_toggle #(.COVER_INDEX(3920)) toggle_3920 (
    .clock(toggle_3920_clock),
    .reset(toggle_3920_reset),
    .valid(toggle_3920_valid)
  );
  assign io_in_ready = state == 3'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 129:25]
  assign io_out_valid = state == 3'h4; // @[src/main/scala/nutcore/backend/fu/MDU.scala 128:39]
  assign io_out_bits = {resR,resQ}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 126:21]
  assign toggle_3657_clock = clock;
  assign toggle_3657_reset = reset;
  assign toggle_3657_valid = state ^ toggle_3657_valid_reg;
  assign toggle_3660_clock = clock;
  assign toggle_3660_reset = reset;
  assign toggle_3660_valid = shiftReg ^ toggle_3660_valid_reg;
  assign toggle_3789_clock = clock;
  assign toggle_3789_reset = reset;
  assign toggle_3789_valid = aSignReg ^ toggle_3789_valid_reg;
  assign toggle_3790_clock = clock;
  assign toggle_3790_reset = reset;
  assign toggle_3790_valid = qSignReg ^ toggle_3790_valid_reg;
  assign toggle_3791_clock = clock;
  assign toggle_3791_reset = reset;
  assign toggle_3791_valid = bReg ^ toggle_3791_valid_reg;
  assign toggle_3855_clock = clock;
  assign toggle_3855_reset = reset;
  assign toggle_3855_valid = aValx2Reg ^ toggle_3855_valid_reg;
  assign toggle_3920_clock = clock;
  assign toggle_3920_reset = reset;
  assign toggle_3920_valid = cnt_value ^ toggle_3920_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
      state <= 3'h0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
    end else if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 95:17]
      state <= 3'h1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 96:11]
    end else if (state == 3'h1) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 97:34]
      state <= 3'h2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 110:11]
    end else if (state == 3'h2) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 111:35]
      state <= 3'h3; // @[src/main/scala/nutcore/backend/fu/MDU.scala 113:11]
    end else begin
      state <= _GEN_8;
    end
    if (!(newReq)) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 95:17]
      if (!(state == 3'h1)) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 97:34]
        if (state == 3'h2) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 111:35]
          shiftReg <= {{1'd0}, _shiftReg_T}; // @[src/main/scala/nutcore/backend/fu/MDU.scala 112:14]
        end else if (state == 3'h3) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 114:37]
          shiftReg <= _shiftReg_T_5; // @[src/main/scala/nutcore/backend/fu/MDU.scala 116:14]
        end
      end
    end
    if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 89:27]
      aSignReg <= aSign; // @[src/main/scala/nutcore/backend/fu/MDU.scala 89:27]
    end
    if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 90:27]
      qSignReg <= (aSign ^ bSign) & ~divBy0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 90:27]
    end
    if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
      if (bSign) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 73:12]
        bReg <= _T_3;
      end else begin
        bReg <= io_in_bits_1;
      end
    end
    if (newReq) begin // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
      aValx2Reg <= _aValx2Reg_T; // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    cnt_value <= _GEN_23[5:0]; // @[src/main/scala/chisel3/util/Counter.scala 61:{40,40}]
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    state_p <= state; // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
    toggle_3657_valid_reg <= state;
    shiftReg_p <= shiftReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    toggle_3660_valid_reg <= shiftReg;
    aSignReg_p <= aSignReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 89:27]
    toggle_3789_valid_reg <= aSignReg;
    qSignReg_p <= qSignReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 90:27]
    toggle_3790_valid_reg <= qSignReg;
    bReg_p <= bReg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    toggle_3791_valid_reg <= bReg;
    aValx2Reg_p <= aValx2Reg; // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    toggle_3855_valid_reg <= aValx2Reg;
    cnt_value_p <= cnt_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    toggle_3920_valid_reg <= cnt_value;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {5{`RANDOM}};
  shiftReg = _RAND_1[128:0];
  _RAND_2 = {1{`RANDOM}};
  aSignReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  qSignReg = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  bReg = _RAND_4[63:0];
  _RAND_5 = {3{`RANDOM}};
  aValx2Reg = _RAND_5[64:0];
  _RAND_6 = {1{`RANDOM}};
  cnt_value = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  state_p = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  toggle_3657_valid_reg = _RAND_8[2:0];
  _RAND_9 = {5{`RANDOM}};
  shiftReg_p = _RAND_9[128:0];
  _RAND_10 = {5{`RANDOM}};
  toggle_3660_valid_reg = _RAND_10[128:0];
  _RAND_11 = {1{`RANDOM}};
  aSignReg_p = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  toggle_3789_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  qSignReg_p = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  toggle_3790_valid_reg = _RAND_14[0:0];
  _RAND_15 = {2{`RANDOM}};
  bReg_p = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  toggle_3791_valid_reg = _RAND_16[63:0];
  _RAND_17 = {3{`RANDOM}};
  aValx2Reg_p = _RAND_17[64:0];
  _RAND_18 = {3{`RANDOM}};
  toggle_3855_valid_reg = _RAND_18[64:0];
  _RAND_19 = {1{`RANDOM}};
  cnt_value_p = _RAND_19[5:0];
  _RAND_20 = {1{`RANDOM}};
  toggle_3920_valid_reg = _RAND_20[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(state_t[0]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[1]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[2]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 77:22]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[0]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[1]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[2]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[3]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[4]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[5]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[6]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[7]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[8]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[9]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[10]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[11]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[12]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[13]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[14]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[15]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[16]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[17]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[18]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[19]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[20]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[21]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[22]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[23]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[24]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[25]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[26]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[27]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[28]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[29]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[30]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[31]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[32]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[33]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[34]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[35]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[36]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[37]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[38]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[39]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[40]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[41]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[42]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[43]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[44]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[45]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[46]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[47]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[48]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[49]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[50]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[51]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[52]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[53]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[54]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[55]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[56]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[57]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[58]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[59]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[60]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[61]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[62]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[63]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[64]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[65]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[66]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[67]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[68]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[69]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[70]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[71]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[72]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[73]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[74]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[75]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[76]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[77]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[78]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[79]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[80]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[81]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[82]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[83]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[84]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[85]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[86]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[87]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[88]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[89]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[90]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[91]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[92]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[93]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[94]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[95]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[96]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[97]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[98]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[99]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[100]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[101]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[102]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[103]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[104]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[105]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[106]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[107]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[108]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[109]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[110]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[111]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[112]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[113]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[114]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[115]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[116]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[117]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[118]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[119]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[120]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[121]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[122]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[123]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[124]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[125]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[126]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[127]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(shiftReg_t[128]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 83:21]
    end
    //
    if (enToggle_past) begin
      cover(aSignReg_t); // @[src/main/scala/nutcore/backend/fu/MDU.scala 89:27]
    end
    //
    if (enToggle_past) begin
      cover(qSignReg_t); // @[src/main/scala/nutcore/backend/fu/MDU.scala 90:27]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[0]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[1]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[2]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[3]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[4]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[5]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[6]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[7]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[8]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[9]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[10]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[11]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[12]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[13]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[14]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[15]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[16]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[17]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[18]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[19]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[20]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[21]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[22]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[23]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[24]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[25]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[26]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[27]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[28]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[29]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[30]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[31]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[32]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[33]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[34]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[35]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[36]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[37]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[38]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[39]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[40]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[41]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[42]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[43]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[44]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[45]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[46]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[47]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[48]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[49]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[50]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[51]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[52]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[53]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[54]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[55]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[56]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[57]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[58]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[59]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[60]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[61]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[62]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(bReg_t[63]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 91:23]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[0]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[1]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[2]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[3]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[4]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[5]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[6]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[7]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[8]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[9]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[10]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[11]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[12]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[13]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[14]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[15]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[16]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[17]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[18]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[19]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[20]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[21]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[22]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[23]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[24]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[25]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[26]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[27]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[28]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[29]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[30]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[31]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[32]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[33]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[34]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[35]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[36]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[37]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[38]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[39]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[40]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[41]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[42]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[43]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[44]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[45]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[46]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[47]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[48]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[49]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[50]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[51]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[52]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[53]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[54]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[55]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[56]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[57]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[58]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[59]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[60]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[61]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[62]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[63]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(aValx2Reg_t[64]); // @[src/main/scala/nutcore/backend/fu/MDU.scala 92:28]
    end
    //
    if (enToggle_past) begin
      cover(cnt_value_t[0]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(cnt_value_t[1]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(cnt_value_t[2]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(cnt_value_t[3]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(cnt_value_t[4]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(cnt_value_t[5]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
  end
endmodule
module MDU(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input         io_in_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input  [63:0] io_in_bits_src1, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input  [63:0] io_in_bits_src2, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input  [6:0]  io_in_bits_func, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
  output [63:0] io_out_bits // @[src/main/scala/nutcore/backend/fu/MDU.scala 136:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  mul_clock; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_reset; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_io_in_ready; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_io_in_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire [64:0] mul_io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire [64:0] mul_io_in_bits_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_io_out_ready; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  mul_io_out_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire [129:0] mul_io_out_bits; // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
  wire  div_clock; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_reset; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_io_in_ready; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_io_in_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire [63:0] div_io_in_bits_0; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire [63:0] div_io_in_bits_1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_io_sign; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  div_io_out_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire [127:0] div_io_out_bits; // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
  wire  isDiv = io_in_bits_func[2]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 41:27]
  wire  isDivSign = isDiv & ~io_in_bits_func[0]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 42:39]
  wire  isW = io_in_bits_func[3]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 43:25]
  wire [64:0] _mul_io_in_bits_0_T_1 = {1'h0,io_in_bits_src1}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  mul_io_in_bits_0_signBit = io_in_bits_src1[63]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [64:0] _mul_io_in_bits_0_T_2 = {mul_io_in_bits_0_signBit,io_in_bits_src1}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  _mul_io_in_bits_0_T_5 = 2'h0 == io_in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _mul_io_in_bits_0_T_6 = 2'h1 == io_in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _mul_io_in_bits_0_T_7 = 2'h2 == io_in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _mul_io_in_bits_0_T_8 = 2'h3 == io_in_bits_func[1:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [64:0] _mul_io_in_bits_0_T_9 = _mul_io_in_bits_0_T_5 ? _mul_io_in_bits_0_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_10 = _mul_io_in_bits_0_T_6 ? _mul_io_in_bits_0_T_2 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_11 = _mul_io_in_bits_0_T_7 ? _mul_io_in_bits_0_T_2 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_12 = _mul_io_in_bits_0_T_8 ? _mul_io_in_bits_0_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_13 = _mul_io_in_bits_0_T_9 | _mul_io_in_bits_0_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_0_T_14 = _mul_io_in_bits_0_T_13 | _mul_io_in_bits_0_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_1 = {1'h0,io_in_bits_src2}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  mul_io_in_bits_1_signBit = io_in_bits_src2[63]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [64:0] _mul_io_in_bits_1_T_2 = {mul_io_in_bits_1_signBit,io_in_bits_src2}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [64:0] _mul_io_in_bits_1_T_9 = _mul_io_in_bits_0_T_5 ? _mul_io_in_bits_1_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_10 = _mul_io_in_bits_0_T_6 ? _mul_io_in_bits_1_T_2 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_11 = _mul_io_in_bits_0_T_7 ? _mul_io_in_bits_1_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_12 = _mul_io_in_bits_0_T_8 ? _mul_io_in_bits_1_T_1 : 65'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_13 = _mul_io_in_bits_1_T_9 | _mul_io_in_bits_1_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [64:0] _mul_io_in_bits_1_T_14 = _mul_io_in_bits_1_T_13 | _mul_io_in_bits_1_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  div_io_in_bits_0_signBit = io_in_bits_src1[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _div_io_in_bits_0_T_1 = div_io_in_bits_0_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _div_io_in_bits_0_T_2 = {_div_io_in_bits_0_T_1,io_in_bits_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _div_io_in_bits_0_T_4 = {32'h0,io_in_bits_src1[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _div_io_in_bits_0_T_5 = isDivSign ? _div_io_in_bits_0_T_2 : _div_io_in_bits_0_T_4; // @[src/main/scala/nutcore/backend/fu/MDU.scala 169:47]
  wire  div_io_in_bits_1_signBit = io_in_bits_src2[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _div_io_in_bits_1_T_1 = div_io_in_bits_1_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _div_io_in_bits_1_T_2 = {_div_io_in_bits_1_T_1,io_in_bits_src2[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _div_io_in_bits_1_T_4 = {32'h0,io_in_bits_src2[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _div_io_in_bits_1_T_5 = isDivSign ? _div_io_in_bits_1_T_2 : _div_io_in_bits_1_T_4; // @[src/main/scala/nutcore/backend/fu/MDU.scala 169:47]
  wire [63:0] mulRes = io_in_bits_func[1:0] == 2'h0 ? mul_io_out_bits[63:0] : mul_io_out_bits[127:64]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 176:19]
  wire [63:0] divRes = io_in_bits_func[1] ? div_io_out_bits[127:64] : div_io_out_bits[63:0]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 177:19]
  wire [63:0] res = isDiv ? divRes : mulRes; // @[src/main/scala/nutcore/backend/fu/MDU.scala 178:16]
  wire  io_out_bits_signBit = res[31]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [31:0] _io_out_bits_T_1 = io_out_bits_signBit ? 32'hffffffff : 32'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _io_out_bits_T_2 = {_io_out_bits_T_1,res[31:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  _isDivReg_T = io_in_ready & io_in_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  isDivReg_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 181:50]
  wire  isDivReg = _isDivReg_T ? isDiv : isDivReg_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 181:21]
  wire  _T = mul_io_out_ready & mul_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  isDivReg_REG_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 181:50]
  wire  isDivReg_REG_t = isDivReg_REG ^ isDivReg_REG_p; // @[src/main/scala/nutcore/backend/fu/MDU.scala 181:50]
  wire  toggle_3926_clock;
  wire  toggle_3926_reset;
  wire  toggle_3926_valid;
  reg  toggle_3926_valid_reg;
  Multiplier mul ( // @[src/main/scala/nutcore/backend/fu/MDU.scala 151:19]
    .clock(mul_clock),
    .reset(mul_reset),
    .io_in_ready(mul_io_in_ready),
    .io_in_valid(mul_io_in_valid),
    .io_in_bits_0(mul_io_in_bits_0),
    .io_in_bits_1(mul_io_in_bits_1),
    .io_out_ready(mul_io_out_ready),
    .io_out_valid(mul_io_out_valid),
    .io_out_bits(mul_io_out_bits)
  );
  Divider div ( // @[src/main/scala/nutcore/backend/fu/MDU.scala 152:19]
    .clock(div_clock),
    .reset(div_reset),
    .io_in_ready(div_io_in_ready),
    .io_in_valid(div_io_in_valid),
    .io_in_bits_0(div_io_in_bits_0),
    .io_in_bits_1(div_io_in_bits_1),
    .io_sign(div_io_sign),
    .io_out_valid(div_io_out_valid),
    .io_out_bits(div_io_out_bits)
  );
  GEN_w1_toggle #(.COVER_INDEX(3926)) toggle_3926 (
    .clock(toggle_3926_clock),
    .reset(toggle_3926_reset),
    .valid(toggle_3926_valid)
  );
  assign io_in_ready = isDiv ? div_io_in_ready : mul_io_in_ready; // @[src/main/scala/nutcore/backend/fu/MDU.scala 182:21]
  assign io_out_valid = isDivReg ? div_io_out_valid : mul_io_out_valid; // @[src/main/scala/nutcore/backend/fu/MDU.scala 183:22]
  assign io_out_bits = isW ? _io_out_bits_T_2 : res; // @[src/main/scala/nutcore/backend/fu/MDU.scala 179:21]
  assign mul_clock = clock;
  assign mul_reset = reset;
  assign mul_io_in_valid = io_in_valid & ~isDiv; // @[src/main/scala/nutcore/backend/fu/MDU.scala 173:34]
  assign mul_io_in_bits_0 = _mul_io_in_bits_0_T_14 | _mul_io_in_bits_0_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign mul_io_in_bits_1 = _mul_io_in_bits_1_T_14 | _mul_io_in_bits_1_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign mul_io_out_ready = 1'h1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 155:17]
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_in_valid = io_in_valid & isDiv; // @[src/main/scala/nutcore/backend/fu/MDU.scala 174:34]
  assign div_io_in_bits_0 = isW ? _div_io_in_bits_0_T_5 : io_in_bits_src1; // @[src/main/scala/nutcore/backend/fu/MDU.scala 169:38]
  assign div_io_in_bits_1 = isW ? _div_io_in_bits_1_T_5 : io_in_bits_src2; // @[src/main/scala/nutcore/backend/fu/MDU.scala 169:38]
  assign div_io_sign = isDiv & ~io_in_bits_func[0]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 42:39]
  assign toggle_3926_clock = clock;
  assign toggle_3926_reset = reset;
  assign toggle_3926_valid = isDivReg_REG ^ toggle_3926_valid_reg;
  always @(posedge clock) begin
    isDivReg_REG <= io_in_bits_func[2]; // @[src/main/scala/nutcore/backend/fu/MDU.scala 41:27]
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    isDivReg_REG_p <= isDivReg_REG; // @[src/main/scala/nutcore/backend/fu/MDU.scala 181:50]
    toggle_3926_valid_reg <= isDivReg_REG;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isDivReg_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  isDivReg_REG_p = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  toggle_3926_valid_reg = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(isDivReg_REG_t); // @[src/main/scala/nutcore/backend/fu/MDU.scala 181:50]
    end
  end
endmodule
module DummyDPICWrapper_1(
  input         clock,
  input         reset,
  input  [63:0] io_bits_privilegeMode, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mstatus, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_sstatus, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mepc, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_sepc, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mtval, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_stval, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mtvec, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_stvec, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mcause, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_scause, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_satp, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mip, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mie, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mscratch, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_sscratch, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_mideleg, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_medeleg // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_privilegeMode; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mstatus; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_sstatus; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mepc; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_sepc; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mtval; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_stval; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mtvec; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_stvec; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mcause; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_scause; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_satp; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mip; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mie; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mscratch; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_sscratch; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_mideleg; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_medeleg; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestCSRState dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_privilegeMode(dpic_io_privilegeMode),
    .io_mstatus(dpic_io_mstatus),
    .io_sstatus(dpic_io_sstatus),
    .io_mepc(dpic_io_mepc),
    .io_sepc(dpic_io_sepc),
    .io_mtval(dpic_io_mtval),
    .io_stval(dpic_io_stval),
    .io_mtvec(dpic_io_mtvec),
    .io_stvec(dpic_io_stvec),
    .io_mcause(dpic_io_mcause),
    .io_scause(dpic_io_scause),
    .io_satp(dpic_io_satp),
    .io_mip(dpic_io_mip),
    .io_mie(dpic_io_mie),
    .io_mscratch(dpic_io_mscratch),
    .io_sscratch(dpic_io_sscratch),
    .io_mideleg(dpic_io_mideleg),
    .io_medeleg(dpic_io_medeleg),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = 1'h1; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_privilegeMode = io_bits_privilegeMode; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mstatus = io_bits_mstatus; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_sstatus = io_bits_sstatus; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mepc = io_bits_mepc; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_sepc = io_bits_sepc; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mtval = io_bits_mtval; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_stval = io_bits_stval; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mtvec = io_bits_mtvec; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_stvec = io_bits_stvec; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mcause = io_bits_mcause; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_scause = io_bits_scause; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_satp = io_bits_satp; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mip = io_bits_mip; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mie = io_bits_mie; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mscratch = io_bits_mscratch; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_sscratch = io_bits_sscratch; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_mideleg = io_bits_mideleg; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_medeleg = io_bits_medeleg; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module DummyDPICWrapper_2(
  input         clock,
  input         reset,
  input         io_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [31:0] io_bits_interrupt, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [31:0] io_bits_exception, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_exceptionPC, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [31:0] io_bits_exceptionInst // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_valid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [31:0] dpic_io_interrupt; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [31:0] dpic_io_exception; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_exceptionPC; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [31:0] dpic_io_exceptionInst; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestArchEvent dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_valid(dpic_io_valid),
    .io_interrupt(dpic_io_interrupt),
    .io_exception(dpic_io_exception),
    .io_exceptionPC(dpic_io_exceptionPC),
    .io_exceptionInst(dpic_io_exceptionInst),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = io_valid; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_valid = io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_interrupt = io_bits_interrupt; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_exception = io_bits_exception; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_exceptionPC = io_bits_exceptionPC; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_exceptionInst = io_bits_exceptionInst; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module CSRDiffWrapper(
  input         clock,
  input         reset,
  input  [63:0] io_csrState_privilegeMode, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_mstatus, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_sstatus, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_mepc, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_sepc, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_mtval, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_stval, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_mtvec, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_stvec, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_mcause, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_scause, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_satp, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_mip, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_mie, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_mscratch, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_sscratch, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_mideleg, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_csrState_medeleg, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input         io_archEvent_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [31:0] io_archEvent_interrupt, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [31:0] io_archEvent_exception, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [63:0] io_archEvent_exceptionPC, // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
  input  [31:0] io_archEvent_exceptionInst // @[src/main/scala/nutcore/backend/fu/CSR.scala 1042:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
`endif // RANDOMIZE_REG_INIT
  wire  difftest_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_privilegeMode; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mstatus; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_sstatus; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mepc; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_sepc; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mtval; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_stval; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mtvec; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_stvec; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mcause; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_scause; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_satp; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mip; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mie; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mscratch; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_sscratch; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_mideleg; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_medeleg; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftestArchEvent_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftestArchEvent_module_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftestArchEvent_module_io_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftestArchEvent_module_io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [31:0] difftestArchEvent_module_io_bits_interrupt; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [31:0] difftestArchEvent_module_io_bits_exception; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftestArchEvent_module_io_bits_exceptionPC; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [31:0] difftestArchEvent_module_io_bits_exceptionInst; // @[difftest/src/main/scala/DPIC.scala 299:24]
  reg [63:0] difftest_REG_privilegeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_sstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_stvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_satp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_mip; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_mie; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_mscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_sscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg [63:0] difftest_REG_medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
  reg  difftestArchEvent_REG_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:43]
  reg [31:0] difftestArchEvent_REG_interrupt; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:43]
  reg [31:0] difftestArchEvent_REG_exception; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:43]
  reg [63:0] difftestArchEvent_REG_exceptionPC; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:43]
  reg [31:0] difftestArchEvent_REG_exceptionInst; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:43]
  reg  difftestArchEvent_REG_1_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:35]
  reg [31:0] difftestArchEvent_REG_1_interrupt; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:35]
  reg [31:0] difftestArchEvent_REG_1_exception; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:35]
  reg [63:0] difftestArchEvent_REG_1_exceptionPC; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:35]
  reg [31:0] difftestArchEvent_REG_1_exceptionInst; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:35]
  DummyDPICWrapper_1 difftest_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_clock),
    .reset(difftest_module_reset),
    .io_bits_privilegeMode(difftest_module_io_bits_privilegeMode),
    .io_bits_mstatus(difftest_module_io_bits_mstatus),
    .io_bits_sstatus(difftest_module_io_bits_sstatus),
    .io_bits_mepc(difftest_module_io_bits_mepc),
    .io_bits_sepc(difftest_module_io_bits_sepc),
    .io_bits_mtval(difftest_module_io_bits_mtval),
    .io_bits_stval(difftest_module_io_bits_stval),
    .io_bits_mtvec(difftest_module_io_bits_mtvec),
    .io_bits_stvec(difftest_module_io_bits_stvec),
    .io_bits_mcause(difftest_module_io_bits_mcause),
    .io_bits_scause(difftest_module_io_bits_scause),
    .io_bits_satp(difftest_module_io_bits_satp),
    .io_bits_mip(difftest_module_io_bits_mip),
    .io_bits_mie(difftest_module_io_bits_mie),
    .io_bits_mscratch(difftest_module_io_bits_mscratch),
    .io_bits_sscratch(difftest_module_io_bits_sscratch),
    .io_bits_mideleg(difftest_module_io_bits_mideleg),
    .io_bits_medeleg(difftest_module_io_bits_medeleg)
  );
  DummyDPICWrapper_2 difftestArchEvent_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftestArchEvent_module_clock),
    .reset(difftestArchEvent_module_reset),
    .io_valid(difftestArchEvent_module_io_valid),
    .io_bits_valid(difftestArchEvent_module_io_bits_valid),
    .io_bits_interrupt(difftestArchEvent_module_io_bits_interrupt),
    .io_bits_exception(difftestArchEvent_module_io_bits_exception),
    .io_bits_exceptionPC(difftestArchEvent_module_io_bits_exceptionPC),
    .io_bits_exceptionInst(difftestArchEvent_module_io_bits_exceptionInst)
  );
  assign difftest_module_clock = clock;
  assign difftest_module_reset = reset;
  assign difftest_module_io_bits_privilegeMode = difftest_REG_privilegeMode; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_mstatus = difftest_REG_mstatus; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_sstatus = difftest_REG_sstatus; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_mepc = difftest_REG_mepc; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_sepc = difftest_REG_sepc; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_mtval = difftest_REG_mtval; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_stval = difftest_REG_stval; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_mtvec = difftest_REG_mtvec; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_stvec = difftest_REG_stvec; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_mcause = difftest_REG_mcause; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_scause = difftest_REG_scause; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_satp = difftest_REG_satp; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_mip = difftest_REG_mip; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_mie = difftest_REG_mie; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_mscratch = difftest_REG_mscratch; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_sscratch = difftest_REG_sscratch; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_mideleg = difftest_REG_mideleg; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftest_module_io_bits_medeleg = difftest_REG_medeleg; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1048:16]
  assign difftestArchEvent_module_clock = clock;
  assign difftestArchEvent_module_reset = reset;
  assign difftestArchEvent_module_io_valid = difftestArchEvent_REG_1_valid; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1052:25]
  assign difftestArchEvent_module_io_bits_valid = difftestArchEvent_REG_1_valid; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1052:25]
  assign difftestArchEvent_module_io_bits_interrupt = difftestArchEvent_REG_1_interrupt; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1052:25]
  assign difftestArchEvent_module_io_bits_exception = difftestArchEvent_REG_1_exception; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1052:25]
  assign difftestArchEvent_module_io_bits_exceptionPC = difftestArchEvent_REG_1_exceptionPC; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1052:25]
  assign difftestArchEvent_module_io_bits_exceptionInst = difftestArchEvent_REG_1_exceptionInst; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/fu/CSR.scala 1052:25]
  always @(posedge clock) begin
    difftest_REG_privilegeMode <= io_csrState_privilegeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_mstatus <= io_csrState_mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_sstatus <= io_csrState_sstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_mepc <= io_csrState_mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_sepc <= io_csrState_sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_mtval <= io_csrState_mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_stval <= io_csrState_stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_mtvec <= io_csrState_mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_stvec <= io_csrState_stvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_mcause <= io_csrState_mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_scause <= io_csrState_scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_satp <= io_csrState_satp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_mip <= io_csrState_mip; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_mie <= io_csrState_mie; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_mscratch <= io_csrState_mscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_sscratch <= io_csrState_sscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_mideleg <= io_csrState_mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftest_REG_medeleg <= io_csrState_medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1048:26]
    difftestArchEvent_REG_valid <= io_archEvent_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:43]
    difftestArchEvent_REG_interrupt <= io_archEvent_interrupt; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:43]
    difftestArchEvent_REG_exception <= io_archEvent_exception; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:43]
    difftestArchEvent_REG_exceptionPC <= io_archEvent_exceptionPC; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:43]
    difftestArchEvent_REG_exceptionInst <= io_archEvent_exceptionInst; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:43]
    difftestArchEvent_REG_1_valid <= difftestArchEvent_REG_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:35]
    difftestArchEvent_REG_1_interrupt <= difftestArchEvent_REG_interrupt; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:35]
    difftestArchEvent_REG_1_exception <= difftestArchEvent_REG_exception; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:35]
    difftestArchEvent_REG_1_exceptionPC <= difftestArchEvent_REG_exceptionPC; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:35]
    difftestArchEvent_REG_1_exceptionInst <= difftestArchEvent_REG_exceptionInst; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1052:35]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  difftest_REG_privilegeMode = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  difftest_REG_mstatus = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  difftest_REG_sstatus = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  difftest_REG_mepc = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  difftest_REG_sepc = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  difftest_REG_mtval = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  difftest_REG_stval = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  difftest_REG_mtvec = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  difftest_REG_stvec = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  difftest_REG_mcause = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  difftest_REG_scause = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  difftest_REG_satp = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  difftest_REG_mip = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  difftest_REG_mie = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  difftest_REG_mscratch = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  difftest_REG_sscratch = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  difftest_REG_mideleg = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  difftest_REG_medeleg = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  difftestArchEvent_REG_valid = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  difftestArchEvent_REG_interrupt = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  difftestArchEvent_REG_exception = _RAND_20[31:0];
  _RAND_21 = {2{`RANDOM}};
  difftestArchEvent_REG_exceptionPC = _RAND_21[63:0];
  _RAND_22 = {1{`RANDOM}};
  difftestArchEvent_REG_exceptionInst = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  difftestArchEvent_REG_1_valid = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  difftestArchEvent_REG_1_interrupt = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  difftestArchEvent_REG_1_exception = _RAND_25[31:0];
  _RAND_26 = {2{`RANDOM}};
  difftestArchEvent_REG_1_exceptionPC = _RAND_26[63:0];
  _RAND_27 = {1{`RANDOM}};
  difftestArchEvent_REG_1_exceptionInst = _RAND_27[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CSR(
  input         clock,
  input         reset,
  input         io_in_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [63:0] io_in_bits_src1, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [63:0] io_in_bits_src2, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [6:0]  io_in_bits_func, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_out_ready, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_out_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output [63:0] io_out_bits, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [63:0] io_cfIn_instr, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [38:0] io_cfIn_pc, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_1, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_2, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_4, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_5, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_6, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_7, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_12, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_13, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_exceptionVec_15, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_intrVec_1, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_intrVec_3, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_intrVec_5, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_intrVec_7, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_intrVec_9, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_intrVec_11, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_cfIn_crossBoundaryFault, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output [38:0] io_redirect_target, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_redirect_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_instrValid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_illegalJump_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [63:0] io_illegalJump_bits, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input  [63:0] io_dmemExceptionAddr, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_xretIsIllegal_ready, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_xretIsIllegal_valid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output [63:0] io_xretIsIllegal_bits, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output [1:0]  io_imemMMU_priviledgeMode, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output [1:0]  io_dmemMMU_priviledgeMode, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_dmemMMU_status_sum, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_dmemMMU_status_mxr, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_dmemMMU_loadPF, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_dmemMMU_storePF, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_dmemMMU_laf, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_dmemMMU_saf, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_wenFix, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_isPerfRead, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_isExit, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_vmEnable, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         io_rfWenReal, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_sfence_vma_invalid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  output        io_wfi_invalid, // @[src/main/scala/nutcore/backend/fu/CSR.scala 200:14]
  input         set_lr,
  output        lr_0,
  input         meip_0,
  output [63:0] lrAddr_0,
  output [63:0] satp_0,
  input         mtip_0,
  input         perfCntCondMultiCommit,
  input         set_lr_val,
  output [11:0] intrVecIDU_0,
  input  [63:0] set_lr_addr,
  input         msip_0,
  input         perfCntCondMinstret
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
`endif // RANDOMIZE_REG_INIT
  wire  CSRDiffWrapper_clock; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire  CSRDiffWrapper_reset; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_privilegeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_sstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_stvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_satp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mip; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mie; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_sscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_csrState_medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire  CSRDiffWrapper_io_archEvent_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [31:0] CSRDiffWrapper_io_archEvent_interrupt; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [31:0] CSRDiffWrapper_io_archEvent_exception; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [63:0] CSRDiffWrapper_io_archEvent_exceptionPC; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  wire [31:0] CSRDiffWrapper_io_archEvent_exceptionInst; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
  reg [1:0] priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:31]
  reg [63:0] mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
  reg [63:0] mcounteren; // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
  reg [63:0] mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
  reg [63:0] mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
  reg [63:0] mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
  reg [63:0] mie; // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
  reg [63:0] mipReg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
  wire [11:0] _mip_T = {meip_0,1'h0,1'h0,1'h0,mtip_0,1'h0,2'h0,msip_0,3'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:22]
  wire [63:0] _GEN_98 = {{52'd0}, _mip_T}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:29]
  wire [63:0] _mip_T_1 = _GEN_98 | mipReg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:29]
  wire  mip_s_u = _mip_T_1[0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_s_s = _mip_T_1[1]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_s_h = _mip_T_1[2]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_s_m = _mip_T_1[3]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_t_u = _mip_T_1[4]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_t_s = _mip_T_1[5]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_t_h = _mip_T_1[6]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_t_m = _mip_T_1[7]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_e_u = _mip_T_1[8]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_e_s = _mip_T_1[9]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_e_h = _mip_T_1[10]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  wire  mip_e_m = _mip_T_1[11]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 281:47]
  reg [63:0] mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
  wire  mstatusStruct_ie_u = mstatus[0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_ie_s = mstatus[1]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_ie_h = mstatus[2]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_ie_m = mstatus[3]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_pie_u = mstatus[4]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_pie_s = mstatus[5]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_pie_h = mstatus[6]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_pie_m = mstatus[7]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_spp = mstatus[8]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire [1:0] mstatusStruct_hpp = mstatus[10:9]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire [1:0] mstatusStruct_mpp = mstatus[12:11]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire [1:0] mstatusStruct_fs = mstatus[14:13]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire [1:0] mstatusStruct_xs = mstatus[16:15]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_mprv = mstatus[17]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_sum = mstatus[18]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_mxr = mstatus[19]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_tvm = mstatus[20]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_tw = mstatus[21]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_tsr = mstatus[22]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire [8:0] mstatusStruct_pad0 = mstatus[31:23]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire [1:0] mstatusStruct_uxl = mstatus[33:32]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire [1:0] mstatusStruct_sxl = mstatus[35:34]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire [26:0] mstatusStruct_pad1 = mstatus[62:36]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  wire  mstatusStruct_sd = mstatus[63]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  reg [63:0] medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
  reg [63:0] mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
  reg [63:0] mscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
  reg [63:0] stvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
  wire [63:0] sieMask = 64'h222 & mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 379:32]
  reg [63:0] satp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
  wire [3:0] satpStruct_mode = satp[63:60]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 384:33]
  wire  _vmEnable_T_1 = priviledgeMode < 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 251:38]
  wire  vmEnable = satpStruct_mode == 4'h8 & priviledgeMode < 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 251:20]
  reg [63:0] sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
  reg [63:0] scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
  reg [63:0] stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
  reg [63:0] sscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
  reg [63:0] scounteren; // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
  reg  lr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 407:19]
  reg [63:0] lrAddr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
  reg [63:0] perfCnts_0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
  reg [63:0] perfCnts_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
  reg [63:0] perfCnts_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
  wire [5:0] lo = {mip_t_s,mip_t_u,mip_s_m,mip_s_h,mip_s_s,mip_s_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 467:27]
  wire [11:0] _T_25 = {mip_e_m,mip_e_h,mip_e_s,mip_e_u,mip_t_m,mip_t_h,lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 467:27]
  wire [11:0] addr = io_in_bits_src2[11:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 507:18]
  wire [63:0] csri = {59'h0,io_cfIn_instr[19:15]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire  _rdata_T_29 = 12'hf12 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_30 = 12'h180 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_59 = _rdata_T_30 ? satp : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_31 = 12'h140 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_60 = _rdata_T_31 ? sscratch : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_88 = _rdata_T_59 | _rdata_T_60; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_32 = 12'h306 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_61 = _rdata_T_32 ? mcounteren : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_89 = _rdata_T_88 | _rdata_T_61; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_33 = 12'hf11 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_34 = 12'h104 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_5 = mie & sieMask; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_63 = _rdata_T_34 ? _rdata_T_5 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_91 = _rdata_T_89 | _rdata_T_63; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_35 = 12'h144 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _GEN_99 = {{52'd0}, _T_25}; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_6 = _GEN_99 & sieMask; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_64 = _rdata_T_35 ? _rdata_T_6 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_92 = _rdata_T_91 | _rdata_T_64; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_36 = 12'h100 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_7 = mstatus & 64'h80000003000d8122; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_65 = _rdata_T_36 ? _rdata_T_7 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_93 = _rdata_T_92 | _rdata_T_65; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_37 = 12'h305 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_66 = _rdata_T_37 ? mtvec : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_94 = _rdata_T_93 | _rdata_T_66; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_38 = 12'h300 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_9 = mstatus & 64'h8000000f007ff9aa; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_67 = _rdata_T_38 ? _rdata_T_9 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_95 = _rdata_T_94 | _rdata_T_67; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_39 = 12'hf13 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_40 = 12'h340 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_69 = _rdata_T_40 ? mscratch : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_97 = _rdata_T_95 | _rdata_T_69; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_41 = 12'h142 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_70 = _rdata_T_41 ? scause : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_98 = _rdata_T_97 | _rdata_T_70; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_42 = 12'h302 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_71 = _rdata_T_42 ? medeleg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_99 = _rdata_T_98 | _rdata_T_71; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_43 = 12'h105 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_72 = _rdata_T_43 ? stvec : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_100 = _rdata_T_99 | _rdata_T_72; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_44 = 12'h141 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_73 = _rdata_T_44 ? sepc : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_101 = _rdata_T_100 | _rdata_T_73; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_45 = 12'h342 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_74 = _rdata_T_45 ? mcause : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_102 = _rdata_T_101 | _rdata_T_74; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_46 = 12'h304 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_75 = _rdata_T_46 ? mie : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_103 = _rdata_T_102 | _rdata_T_75; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_47 = 12'hb01 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_76 = _rdata_T_47 ? perfCnts_1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_104 = _rdata_T_103 | _rdata_T_76; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_48 = 12'h143 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_77 = _rdata_T_48 ? stval : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_105 = _rdata_T_104 | _rdata_T_77; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_49 = 12'h301 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_78 = _rdata_T_49 ? 64'h8000000000141105 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_106 = _rdata_T_105 | _rdata_T_78; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_50 = 12'hb00 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_79 = _rdata_T_50 ? perfCnts_0 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_107 = _rdata_T_106 | _rdata_T_79; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_51 = 12'h344 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_22 = {{52'd0}, _T_25}; // @[src/main/scala/utils/RegMap.scala 48:84]
  wire [63:0] _rdata_T_80 = _rdata_T_51 ? _rdata_T_22 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_108 = _rdata_T_107 | _rdata_T_80; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_52 = 12'hb02 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_81 = _rdata_T_52 ? perfCnts_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_109 = _rdata_T_108 | _rdata_T_81; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_53 = 12'h303 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_82 = _rdata_T_53 ? mideleg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_110 = _rdata_T_109 | _rdata_T_82; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_54 = 12'hf14 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_55 = 12'h341 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_84 = _rdata_T_55 ? mepc : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_112 = _rdata_T_110 | _rdata_T_84; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_56 = 12'h343 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_85 = _rdata_T_56 ? mtval : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _rdata_T_113 = _rdata_T_112 | _rdata_T_85; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _rdata_T_57 = 12'h106 == addr; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _rdata_T_86 = _rdata_T_57 ? scounteren : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdata = _rdata_T_113 | _rdata_T_86; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T = rdata | io_in_bits_src1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 512:30]
  wire [63:0] _wdata_T_1 = ~io_in_bits_src1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 513:33]
  wire [63:0] _wdata_T_2 = rdata & _wdata_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 513:30]
  wire [63:0] _wdata_T_3 = rdata | csri; // @[src/main/scala/nutcore/backend/fu/CSR.scala 515:30]
  wire [63:0] _wdata_T_4 = ~csri; // @[src/main/scala/nutcore/backend/fu/CSR.scala 516:33]
  wire [63:0] _wdata_T_5 = rdata & _wdata_T_4; // @[src/main/scala/nutcore/backend/fu/CSR.scala 516:30]
  wire  _wdata_T_6 = 7'h1 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_7 = 7'h2 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_8 = 7'h3 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_9 = 7'h5 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_10 = 7'h6 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _wdata_T_11 = 7'h7 == io_in_bits_func; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _wdata_T_12 = _wdata_T_6 ? io_in_bits_src1 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_13 = _wdata_T_7 ? _wdata_T : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_14 = _wdata_T_8 ? _wdata_T_2 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_15 = _wdata_T_9 ? csri : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_16 = _wdata_T_10 ? _wdata_T_3 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_17 = _wdata_T_11 ? _wdata_T_5 : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_18 = _wdata_T_12 | _wdata_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_19 = _wdata_T_18 | _wdata_T_14; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_20 = _wdata_T_19 | _wdata_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _wdata_T_21 = _wdata_T_20 | _wdata_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] wdata = _wdata_T_21 | _wdata_T_17; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  satpLegalMode = wdata[63:60] == 4'h0 | wdata[63:60] == 4'h8; // @[src/main/scala/nutcore/backend/fu/CSR.scala 522:69]
  wire [7:0] wen_lo = {io_cfIn_exceptionVec_7,io_cfIn_exceptionVec_6,io_cfIn_exceptionVec_5,io_cfIn_exceptionVec_4,1'h0,
    io_cfIn_exceptionVec_2,io_cfIn_exceptionVec_1,1'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 525:45]
  wire [15:0] _wen_T = {io_cfIn_exceptionVec_15,1'h0,io_cfIn_exceptionVec_13,io_cfIn_exceptionVec_12,4'h0,wen_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 525:45]
  wire  _wen_T_2 = ~(|_wen_T); // @[src/main/scala/nutcore/backend/fu/CSR.scala 525:23]
  wire  _wen_T_4 = io_in_bits_func != 7'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 525:64]
  wire  wen = io_in_valid & ~(|_wen_T) & io_in_bits_func != 7'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 525:56]
  wire  isIllegalMode = priviledgeMode < addr[9:8]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 526:39]
  wire  isCSRRS = io_in_bits_func == 7'h2 | io_in_bits_func == 7'h6; // @[src/main/scala/nutcore/backend/fu/CSR.scala 531:40]
  wire  isCSRRC = io_in_bits_func == 7'h3 | io_in_bits_func == 7'h7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 532:40]
  wire  noWriteSideEffect = (isCSRRS | isCSRRC) & io_cfIn_instr[19:15] == 5'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 533:48]
  wire  isIllegalWrite = wen & addr[11:10] == 2'h3 & ~noWriteSideEffect; // @[src/main/scala/nutcore/backend/fu/CSR.scala 535:58]
  wire  _tvm_T_1 = priviledgeMode == 2'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 541:57]
  wire  tvm = mstatusStruct_tvm & priviledgeMode == 2'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 541:39]
  wire  _io_sfence_vma_invalid_T = priviledgeMode == 2'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 542:43]
  wire  _isIllegalTVM_T_1 = addr == 12'h180; // @[src/main/scala/nutcore/backend/fu/CSR.scala 543:42]
  wire  isIllegalTVM = tvm & wen & addr == 12'h180; // @[src/main/scala/nutcore/backend/fu/CSR.scala 543:34]
  wire  isIllegalAccess = isIllegalMode | isIllegalWrite | isIllegalTVM; // @[src/main/scala/nutcore/backend/fu/CSR.scala 544:57]
  wire  _canWriteCSR_T = ~isIllegalAccess; // @[src/main/scala/nutcore/backend/fu/CSR.scala 548:28]
  wire  _canWriteCSR_T_1 = wen & ~isIllegalAccess; // @[src/main/scala/nutcore/backend/fu/CSR.scala 548:25]
  wire  canWriteCSR = wen & ~isIllegalAccess & (addr != 12'h180 | satpLegalMode); // @[src/main/scala/nutcore/backend/fu/CSR.scala 548:45]
  wire [63:0] _satp_T = wdata & 64'h8ffff000000fffff; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _satp_T_2 = satp & 64'h70000ffffff00000; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _satp_T_3 = _satp_T | _satp_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _mie_T = wdata & sieMask; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mie_T_1 = ~sieMask; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [63:0] _mie_T_2 = mie & _mie_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mie_T_3 = _mie_T | _mie_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _mstatus_T = wdata & 64'hc0122; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mstatus_T_2 = mstatus & 64'hfffffffffff3fedd; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mstatus_T_3 = _mstatus_T | _mstatus_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [1:0] mstatus_mstatusOld_mpp = _mstatus_T_3[12:11]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 320:47]
  wire [1:0] mstatus_mstatusOld_fs = _mstatus_T_3[14:13]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 320:47]
  wire [1:0] mstatus_mppFix = mstatus_mstatusOld_mpp == 2'h2 ? 2'h0 : mstatus_mstatusOld_mpp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 324:21]
  wire [63:0] mstatus_mstatusNew = {mstatus_mstatusOld_fs == 2'h3,_mstatus_T_3[62:13],mstatus_mppFix,_mstatus_T_3[10:0]}
    ; // @[src/main/scala/nutcore/backend/fu/CSR.scala 325:25]
  wire [63:0] _GEN_6 = canWriteCSR & addr == 12'h100 ? mstatus_mstatusNew : mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _mtvec_T = wdata & 64'hfffffffffffffffc; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mtvec_T_2 = mtvec & 64'h3; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mtvec_T_3 = _mtvec_T | _mtvec_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _mstatus_T_4 = wdata & 64'h80000000007e19aa; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mstatus_T_6 = mstatus & 64'h7fffffffff81e655; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mstatus_T_7 = _mstatus_T_4 | _mstatus_T_6; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [1:0] mstatus_mstatusOld_1_mpp = _mstatus_T_7[12:11]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 320:47]
  wire [1:0] mstatus_mstatusOld_1_fs = _mstatus_T_7[14:13]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 320:47]
  wire [1:0] mstatus_mppFix_1 = mstatus_mstatusOld_1_mpp == 2'h2 ? 2'h0 : mstatus_mstatusOld_1_mpp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 324:21]
  wire [63:0] mstatus_mstatusNew_1 = {mstatus_mstatusOld_1_fs == 2'h3,_mstatus_T_7[62:13],mstatus_mppFix_1,_mstatus_T_7[
    10:0]}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 325:25]
  wire [63:0] _GEN_8 = canWriteCSR & addr == 12'h300 ? mstatus_mstatusNew_1 : _GEN_6; // @[src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _GEN_10 = canWriteCSR & addr == 12'h142 ? wdata : scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire  _T_65 = addr == 12'h302; // @[src/main/scala/utils/RegMap.scala 50:65]
  wire [63:0] _medeleg_T = wdata & 64'hb3ff; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _medeleg_T_2 = medeleg & 64'hffffffffffff4c00; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _medeleg_T_3 = _medeleg_T | _medeleg_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _stvec_T_2 = stvec & 64'h3; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _stvec_T_3 = _mtvec_T | _stvec_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _sepc_T = wdata & 64'hfffffffffffffffe; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _sepc_T_2 = sepc & 64'h1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _sepc_T_3 = _sepc_T | _sepc_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _GEN_13 = canWriteCSR & addr == 12'h141 ? _sepc_T_3 : sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _GEN_14 = canWriteCSR & addr == 12'h342 ? wdata : mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _mie_T_4 = wdata & 64'haaa; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mie_T_6 = mie & 64'hfffffffffffff555; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mie_T_7 = _mie_T_4 | _mie_T_6; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _GEN_17 = canWriteCSR & addr == 12'h143 ? wdata : stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire  _T_79 = addr == 12'hb00; // @[src/main/scala/utils/RegMap.scala 50:65]
  wire  _T_81 = addr == 12'hb02; // @[src/main/scala/utils/RegMap.scala 50:65]
  wire [63:0] _mideleg_T = wdata & 64'h222; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mideleg_T_2 = mideleg & 64'hfffffffffffffddd; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mideleg_T_3 = _mideleg_T | _mideleg_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _mepc_T_2 = mepc & 64'h1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mepc_T_3 = _sepc_T | _mepc_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _GEN_21 = canWriteCSR & addr == 12'h341 ? _mepc_T_3 : mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire [63:0] _GEN_22 = canWriteCSR & addr == 12'h343 ? wdata : mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22 src/main/scala/utils/RegMap.scala 50:{72,76}]
  wire  _isIllegalAddr_illegalAddr_T_1 = _rdata_T_29 ? 1'h0 : 1'h1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_3 = _rdata_T_30 ? 1'h0 : _isIllegalAddr_illegalAddr_T_1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_5 = _rdata_T_31 ? 1'h0 : _isIllegalAddr_illegalAddr_T_3; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_7 = _rdata_T_32 ? 1'h0 : _isIllegalAddr_illegalAddr_T_5; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_9 = _rdata_T_33 ? 1'h0 : _isIllegalAddr_illegalAddr_T_7; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_11 = _rdata_T_34 ? 1'h0 : _isIllegalAddr_illegalAddr_T_9; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_13 = _rdata_T_35 ? 1'h0 : _isIllegalAddr_illegalAddr_T_11; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_15 = _rdata_T_36 ? 1'h0 : _isIllegalAddr_illegalAddr_T_13; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_17 = _rdata_T_37 ? 1'h0 : _isIllegalAddr_illegalAddr_T_15; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_19 = _rdata_T_38 ? 1'h0 : _isIllegalAddr_illegalAddr_T_17; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_21 = _rdata_T_39 ? 1'h0 : _isIllegalAddr_illegalAddr_T_19; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_23 = _rdata_T_40 ? 1'h0 : _isIllegalAddr_illegalAddr_T_21; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_25 = _rdata_T_41 ? 1'h0 : _isIllegalAddr_illegalAddr_T_23; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_27 = _rdata_T_42 ? 1'h0 : _isIllegalAddr_illegalAddr_T_25; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_29 = _rdata_T_43 ? 1'h0 : _isIllegalAddr_illegalAddr_T_27; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_31 = _rdata_T_44 ? 1'h0 : _isIllegalAddr_illegalAddr_T_29; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_33 = _rdata_T_45 ? 1'h0 : _isIllegalAddr_illegalAddr_T_31; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_35 = _rdata_T_46 ? 1'h0 : _isIllegalAddr_illegalAddr_T_33; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_37 = _rdata_T_47 ? 1'h0 : _isIllegalAddr_illegalAddr_T_35; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_39 = _rdata_T_48 ? 1'h0 : _isIllegalAddr_illegalAddr_T_37; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_41 = _rdata_T_49 ? 1'h0 : _isIllegalAddr_illegalAddr_T_39; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_43 = _rdata_T_50 ? 1'h0 : _isIllegalAddr_illegalAddr_T_41; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_45 = _rdata_T_51 ? 1'h0 : _isIllegalAddr_illegalAddr_T_43; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_47 = _rdata_T_52 ? 1'h0 : _isIllegalAddr_illegalAddr_T_45; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_49 = _rdata_T_53 ? 1'h0 : _isIllegalAddr_illegalAddr_T_47; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_51 = _rdata_T_54 ? 1'h0 : _isIllegalAddr_illegalAddr_T_49; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_53 = _rdata_T_55 ? 1'h0 : _isIllegalAddr_illegalAddr_T_51; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _isIllegalAddr_illegalAddr_T_55 = _rdata_T_56 ? 1'h0 : _isIllegalAddr_illegalAddr_T_53; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  isIllegalAddr = _rdata_T_57 ? 1'h0 : _isIllegalAddr_illegalAddr_T_55; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  resetSatp = _isIllegalTVM_T_1 & wen & _canWriteCSR_T; // @[src/main/scala/nutcore/backend/fu/CSR.scala 552:42]
  wire  _io_isExit_T = addr == 12'h344; // @[src/main/scala/nutcore/backend/fu/CSR.scala 555:38]
  wire  _io_isExit_T_1 = addr == 12'h144; // @[src/main/scala/nutcore/backend/fu/CSR.scala 555:56]
  wire  _io_isExit_T_9 = _canWriteCSR_T_1 | ~wen; // @[src/main/scala/nutcore/backend/fu/CSR.scala 556:30]
  wire  _io_isExit_T_10 = io_out_valid & (addr == 12'h344 | addr == 12'h144) & _wen_T_4 & _io_isExit_T_9; // @[src/main/scala/nutcore/backend/fu/CSR.scala 555:93]
  wire [63:0] _mipReg_T = wdata & 64'h77f; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _mipReg_T_2 = mipReg & 64'hfffffffffffff880; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mipReg_T_3 = _mipReg_T | _mipReg_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _mipReg_T_6 = mipReg & _mie_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mipReg_T_7 = _mie_T | _mipReg_T_6; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _isEbreak_T_1 = io_in_bits_func == 7'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 568:46]
  wire  isEbreak = addr == 12'h1 & io_in_bits_func == 7'h0 & _wen_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 568:90]
  wire  isEcall = addr == 12'h0 & _isEbreak_T_1 & _wen_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 569:88]
  wire  isMret = _T_65 & _isEbreak_T_1 & _wen_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 570:88]
  wire  isSret = addr == 12'h102 & _isEbreak_T_1 & _wen_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 571:88]
  wire  isUret = addr == 12'h2 & _isEbreak_T_1 & _wen_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 572:88]
  wire  hasInstrPageFault = io_cfIn_exceptionVec_12 & io_instrValid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 632:63]
  wire  hasInstrAccessFault = io_cfIn_exceptionVec_1 & io_instrValid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 633:67]
  wire  hasLoadPageFault = io_dmemMMU_loadPF | io_cfIn_exceptionVec_13; // @[src/main/scala/nutcore/backend/fu/CSR.scala 634:43]
  wire  hasStorePageFault = io_dmemMMU_storePF | io_cfIn_exceptionVec_15; // @[src/main/scala/nutcore/backend/fu/CSR.scala 635:45]
  wire  hasLoadAccessFault = io_dmemMMU_laf | io_cfIn_exceptionVec_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 636:42]
  wire  hasStoreAccessFault = io_dmemMMU_saf | io_cfIn_exceptionVec_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 637:43]
  wire [38:0] _imemExceptionAddr_T_1 = io_cfIn_pc + 39'h2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 644:42]
  wire  imemExceptionAddr_signBit = _imemExceptionAddr_T_1[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _imemExceptionAddr_T_2 = imemExceptionAddr_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imemExceptionAddr_T_3 = {_imemExceptionAddr_T_2,_imemExceptionAddr_T_1}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _imemExceptionAddr_T_6 = {25'h0,_imemExceptionAddr_T_1}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _imemExceptionAddr_T_7 = vmEnable ? _imemExceptionAddr_T_3 : _imemExceptionAddr_T_6; // @[src/main/scala/nutcore/backend/fu/CSR.scala 644:12]
  wire  imemExceptionAddr_signBit_1 = io_cfIn_pc[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _imemExceptionAddr_T_8 = imemExceptionAddr_signBit_1 ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _imemExceptionAddr_T_9 = {_imemExceptionAddr_T_8,io_cfIn_pc}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire [63:0] _imemExceptionAddr_T_10 = {25'h0,io_cfIn_pc}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [63:0] _imemExceptionAddr_T_11 = vmEnable ? _imemExceptionAddr_T_9 : _imemExceptionAddr_T_10; // @[src/main/scala/nutcore/backend/fu/CSR.scala 645:12]
  wire [63:0] _imemExceptionAddr_T_12 = io_cfIn_crossBoundaryFault ? _imemExceptionAddr_T_7 : _imemExceptionAddr_T_11; // @[src/main/scala/nutcore/backend/fu/CSR.scala 643:10]
  wire [63:0] imemExceptionAddr = io_illegalJump_valid ? io_illegalJump_bits : _imemExceptionAddr_T_12; // @[src/main/scala/nutcore/backend/fu/CSR.scala 641:29]
  wire  mipRaiseIntr_e_s = mip_e_s | meip_0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 672:31]
  wire [11:0] _ideleg_T = {mip_e_m,mip_e_h,mipRaiseIntr_e_s,mip_e_u,mip_t_m,mip_t_h,lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 674:41]
  wire [63:0] _GEN_100 = {{52'd0}, _ideleg_T}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 674:26]
  wire [63:0] ideleg = mideleg & _GEN_100; // @[src/main/scala/nutcore/backend/fu/CSR.scala 674:26]
  wire  _intrVecEnable_0_T_2 = priviledgeMode < 2'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:125]
  wire  _intrVecEnable_0_T_4 = priviledgeMode == 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 676:53]
  wire  _intrVecEnable_0_T_7 = priviledgeMode == 2'h3 & mstatusStruct_ie_m | _vmEnable_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 676:87]
  wire  intrVecEnable_0 = ideleg[0] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_1 = ideleg[1] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_2 = ideleg[2] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_3 = ideleg[3] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_4 = ideleg[4] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_5 = ideleg[5] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_6 = ideleg[6] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_7 = ideleg[7] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_8 = ideleg[8] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_9 = ideleg[9] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_10 = ideleg[10] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire  intrVecEnable_11 = ideleg[11] ? _tvm_T_1 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _intrVecEnable_0_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 675:51]
  wire [11:0] _intrVec_T_2 = mie[11:0] & _ideleg_T; // @[src/main/scala/nutcore/backend/fu/CSR.scala 680:27]
  wire [5:0] intrVec_lo_1 = {intrVecEnable_5,intrVecEnable_4,intrVecEnable_3,intrVecEnable_2,intrVecEnable_1,
    intrVecEnable_0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 680:65]
  wire [11:0] _intrVec_T_3 = {intrVecEnable_11,intrVecEnable_10,intrVecEnable_9,intrVecEnable_8,intrVecEnable_7,
    intrVecEnable_6,intrVec_lo_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 680:65]
  wire [11:0] intrVec = _intrVec_T_2 & _intrVec_T_3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 680:49]
  wire [5:0] intrVecIDU_lo = {intrVec[5],1'h0,intrVec[3],1'h0,intrVec[1],1'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 681:100]
  wire [11:0] intrVecIDU = {intrVec[11],1'h0,intrVec[9],1'h0,intrVec[7],1'h0,intrVecIDU_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 681:100]
  wire [2:0] _intrNO_T = io_cfIn_intrVec_5 ? 3'h5 : 3'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 685:69]
  wire [3:0] _intrNO_T_1 = io_cfIn_intrVec_9 ? 4'h9 : {{1'd0}, _intrNO_T}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 685:69]
  wire [3:0] _intrNO_T_2 = io_cfIn_intrVec_1 ? 4'h1 : _intrNO_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 685:69]
  wire [3:0] _intrNO_T_3 = io_cfIn_intrVec_7 ? 4'h7 : _intrNO_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 685:69]
  wire [3:0] _intrNO_T_4 = io_cfIn_intrVec_11 ? 4'hb : _intrNO_T_3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 685:69]
  wire [3:0] intrNO = io_cfIn_intrVec_3 ? 4'h3 : _intrNO_T_4; // @[src/main/scala/nutcore/backend/fu/CSR.scala 685:69]
  wire [5:0] _raiseIntr_T = {io_cfIn_intrVec_5,io_cfIn_intrVec_9,io_cfIn_intrVec_1,io_cfIn_intrVec_7,io_cfIn_intrVec_11,
    io_cfIn_intrVec_3}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 687:69]
  wire  raiseIntr = |_raiseIntr_T; // @[src/main/scala/nutcore/backend/fu/CSR.scala 687:76]
  wire  _illegalMret_T = io_in_valid & isMret; // @[src/main/scala/nutcore/backend/fu/CSR.scala 690:33]
  wire  illegalMret = io_in_valid & isMret & _vmEnable_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 690:43]
  wire  _illegalSret_T = io_in_valid & isSret; // @[src/main/scala/nutcore/backend/fu/CSR.scala 691:33]
  wire  illegalSret = io_in_valid & isSret & _intrVecEnable_0_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 691:43]
  wire  illegalSModeSret = _illegalSret_T & _tvm_T_1 & mstatusStruct_tsr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 692:76]
  wire  isIllegalPrivOp = illegalMret | illegalSret | illegalSModeSret; // @[src/main/scala/nutcore/backend/fu/CSR.scala 693:52]
  wire  csrExceptionVec_3 = io_in_valid & isEbreak; // @[src/main/scala/nutcore/backend/fu/CSR.scala 698:46]
  wire  csrExceptionVec_11 = _intrVecEnable_0_T_4 & io_in_valid & isEcall; // @[src/main/scala/nutcore/backend/fu/CSR.scala 699:70]
  wire  csrExceptionVec_9 = _tvm_T_1 & io_in_valid & isEcall; // @[src/main/scala/nutcore/backend/fu/CSR.scala 700:70]
  wire  csrExceptionVec_8 = _io_sfence_vma_invalid_T & io_in_valid & isEcall; // @[src/main/scala/nutcore/backend/fu/CSR.scala 701:70]
  wire  csrExceptionVec_2 = (isIllegalAddr | isIllegalAccess) & wen | isIllegalPrivOp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 702:79]
  wire [7:0] raiseExceptionVec_lo = {hasStoreAccessFault,1'h0,hasLoadAccessFault,1'h0,csrExceptionVec_3,
    csrExceptionVec_2,hasInstrAccessFault,1'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 709:43]
  wire [15:0] _raiseExceptionVec_T = {hasStorePageFault,1'h0,hasLoadPageFault,1'h0,csrExceptionVec_11,1'h0,
    csrExceptionVec_9,csrExceptionVec_8,raiseExceptionVec_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 709:43]
  wire [15:0] raiseExceptionVec = _raiseExceptionVec_T | _wen_T; // @[src/main/scala/nutcore/backend/fu/CSR.scala 709:50]
  wire  raiseException = |raiseExceptionVec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 710:42]
  wire [2:0] _exceptionNO_T_1 = raiseExceptionVec[5] ? 3'h5 : 3'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [2:0] _exceptionNO_T_3 = raiseExceptionVec[7] ? 3'h7 : _exceptionNO_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_5 = raiseExceptionVec[13] ? 4'hd : {{1'd0}, _exceptionNO_T_3}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_7 = raiseExceptionVec[15] ? 4'hf : _exceptionNO_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_9 = raiseExceptionVec[4] ? 4'h4 : _exceptionNO_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_11 = raiseExceptionVec[6] ? 4'h6 : _exceptionNO_T_9; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_13 = raiseExceptionVec[8] ? 4'h8 : _exceptionNO_T_11; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_15 = raiseExceptionVec[9] ? 4'h9 : _exceptionNO_T_13; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_17 = raiseExceptionVec[11] ? 4'hb : _exceptionNO_T_15; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_19 = raiseExceptionVec[0] ? 4'h0 : _exceptionNO_T_17; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_21 = raiseExceptionVec[2] ? 4'h2 : _exceptionNO_T_19; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_23 = raiseExceptionVec[1] ? 4'h1 : _exceptionNO_T_21; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] _exceptionNO_T_25 = raiseExceptionVec[12] ? 4'hc : _exceptionNO_T_23; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [3:0] exceptionNO = raiseExceptionVec[3] ? 4'h3 : _exceptionNO_T_25; // @[src/main/scala/nutcore/backend/fu/CSR.scala 711:74]
  wire [63:0] _causeNO_T = {raiseIntr, 63'h0}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 714:28]
  wire [3:0] _causeNO_T_1 = raiseIntr ? intrNO : exceptionNO; // @[src/main/scala/nutcore/backend/fu/CSR.scala 714:53]
  wire [63:0] _GEN_101 = {{60'd0}, _causeNO_T_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 714:48]
  wire [63:0] causeNO = _causeNO_T | _GEN_101; // @[src/main/scala/nutcore/backend/fu/CSR.scala 714:48]
  wire  raiseExceptionIntr = (raiseException | raiseIntr) & io_instrValid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 717:58]
  wire [63:0] _redirectTarget_T_3 = _imemExceptionAddr_T_9 + 64'h4; // @[src/main/scala/nutcore/backend/fu/CSR.scala 721:31]
  wire [63:0] deleg = raiseIntr ? mideleg : medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 758:18]
  wire [63:0] _delegS_T_1 = deleg >> causeNO[3:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 760:21]
  wire  delegS = _delegS_T_1[0] & _vmEnable_T_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 760:36]
  wire [63:0] trapTarget = delegS ? stvec : mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 766:20]
  wire [63:0] _GEN_52 = _illegalSret_T & ~illegalSret & ~illegalSModeSret ? sepc : mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 813:63 826:15]
  wire [63:0] retTarget = io_in_valid & isUret ? 64'h0 : _GEN_52; // @[src/main/scala/nutcore/backend/fu/CSR.scala 829:26 837:15]
  wire [63:0] _redirectTarget_T_4 = raiseExceptionIntr ? trapTarget : retTarget; // @[src/main/scala/nutcore/backend/fu/CSR.scala 722:8]
  wire [63:0] redirectTarget = resetSatp ? _redirectTarget_T_3 : _redirectTarget_T_4; // @[src/main/scala/nutcore/backend/fu/CSR.scala 720:27]
  reg [63:0] redirectTargetReg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
  wire  addrNotLegal_signBit = redirectTargetReg[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _addrNotLegal_T_1 = addrNotLegal_signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire [63:0] _addrNotLegal_T_2 = {_addrNotLegal_T_1,redirectTargetReg[38:0]}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  wire  _addrNotLegal_T_3 = redirectTargetReg != _addrNotLegal_T_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 735:23]
  wire  _addrNotLegal_T_5 = |redirectTargetReg[63:39]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 736:44]
  wire  addrNotLegal = vmEnable ? _addrNotLegal_T_3 : _addrNotLegal_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 734:25]
  reg  hasIllegalXRET; // @[src/main/scala/nutcore/backend/fu/CSR.scala 738:31]
  reg  isIllegalXRET_REG; // @[src/main/scala/nutcore/backend/fu/CSR.scala 739:30]
  wire  isIllegalXRET = isIllegalXRET_REG & addrNotLegal; // @[src/main/scala/nutcore/backend/fu/CSR.scala 739:50]
  wire  _T_162 = io_xretIsIllegal_ready & io_xretIsIllegal_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _GEN_27 = _T_162 ? 1'h0 : hasIllegalXRET; // @[src/main/scala/nutcore/backend/fu/CSR.scala 742:38 743:20 738:31]
  wire  _GEN_28 = isIllegalXRET | _GEN_27; // @[src/main/scala/nutcore/backend/fu/CSR.scala 740:24 741:20]
  wire  isPageFault = hasInstrPageFault | hasLoadPageFault | hasStorePageFault; // @[src/main/scala/nutcore/backend/fu/CSR.scala 761:59]
  wire  isAddrMisAligned = io_cfIn_exceptionVec_4 | io_cfIn_exceptionVec_6; // @[src/main/scala/nutcore/backend/fu/CSR.scala 762:48]
  wire  isAccessFault = hasInstrAccessFault | hasLoadAccessFault | hasStoreAccessFault; // @[src/main/scala/nutcore/backend/fu/CSR.scala 763:65]
  wire [63:0] _GEN_29 = delegS ? io_dmemExceptionAddr : _GEN_17; // @[src/main/scala/nutcore/backend/fu/CSR.scala 771:21 772:15]
  wire [63:0] _GEN_30 = delegS ? _GEN_22 : io_dmemExceptionAddr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 771:21 774:15]
  wire [63:0] tval = hasInstrPageFault ? imemExceptionAddr : io_dmemExceptionAddr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 779:21]
  wire [63:0] _GEN_31 = delegS ? tval : _GEN_17; // @[src/main/scala/nutcore/backend/fu/CSR.scala 780:21 781:15]
  wire [63:0] _GEN_32 = delegS ? _GEN_22 : tval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 780:21 783:15]
  wire [63:0] tval_1 = hasInstrAccessFault ? imemExceptionAddr : io_dmemExceptionAddr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 788:21]
  wire [63:0] _GEN_33 = delegS ? tval_1 : _GEN_17; // @[src/main/scala/nutcore/backend/fu/CSR.scala 789:21 790:15]
  wire [63:0] _GEN_34 = delegS ? _GEN_22 : tval_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 789:21 792:15]
  wire [63:0] _GEN_35 = isAccessFault ? _GEN_33 : _GEN_17; // @[src/main/scala/nutcore/backend/fu/CSR.scala 787:83]
  wire [63:0] _GEN_36 = isAccessFault ? _GEN_34 : _GEN_22; // @[src/main/scala/nutcore/backend/fu/CSR.scala 787:83]
  wire [63:0] _GEN_37 = isPageFault ? _GEN_31 : _GEN_35; // @[src/main/scala/nutcore/backend/fu/CSR.scala 778:77]
  wire [63:0] _GEN_38 = isPageFault ? _GEN_32 : _GEN_36; // @[src/main/scala/nutcore/backend/fu/CSR.scala 778:77]
  wire [63:0] _GEN_39 = isAddrMisAligned ? _GEN_29 : _GEN_37; // @[src/main/scala/nutcore/backend/fu/CSR.scala 770:60]
  wire [63:0] _GEN_40 = isAddrMisAligned ? _GEN_30 : _GEN_38; // @[src/main/scala/nutcore/backend/fu/CSR.scala 770:60]
  wire [63:0] _GEN_41 = io_instrValid ? _GEN_39 : _GEN_17; // @[src/main/scala/nutcore/backend/fu/CSR.scala 769:24]
  wire [63:0] _GEN_42 = io_instrValid ? _GEN_40 : _GEN_22; // @[src/main/scala/nutcore/backend/fu/CSR.scala 769:24]
  wire  mstatusNew_mprv = mstatusStruct_mpp != 2'h3 ? 1'h0 : mstatusStruct_mprv; // @[src/main/scala/nutcore/backend/fu/CSR.scala 803:37 804:23 799:30]
  wire [5:0] mstatus_lo_lo = {mstatusStruct_pie_s,mstatusStruct_pie_u,mstatusStruct_pie_m,mstatusStruct_ie_h,
    mstatusStruct_ie_s,mstatusStruct_ie_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 808:27]
  wire [14:0] mstatus_lo = {mstatusStruct_fs,2'h0,mstatusStruct_hpp,mstatusStruct_spp,1'h1,mstatusStruct_pie_h,
    mstatus_lo_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 808:27]
  wire [6:0] mstatus_hi_lo = {mstatusStruct_tw,mstatusStruct_tvm,mstatusStruct_mxr,mstatusStruct_sum,mstatusNew_mprv,
    mstatusStruct_xs}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 808:27]
  wire [63:0] _mstatus_T_8 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0
    ,mstatusStruct_tsr,mstatus_hi_lo,mstatus_lo}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 808:27]
  wire [1:0] _GEN_44 = _illegalMret_T & ~illegalMret ? mstatusStruct_mpp : priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 797:42 802:20 262:31]
  wire [63:0] _GEN_45 = _illegalMret_T & ~illegalMret ? _mstatus_T_8 : _GEN_8; // @[src/main/scala/nutcore/backend/fu/CSR.scala 797:42 808:13]
  wire [1:0] _priviledgeMode_T = {1'h0,mstatusStruct_spp}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 818:26]
  wire [1:0] _GEN_102 = {{1'd0}, mstatusStruct_spp}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 819:26]
  wire  mstatusNew_1_mprv = _GEN_102 != 2'h3 ? 1'h0 : mstatusStruct_mprv; // @[src/main/scala/nutcore/backend/fu/CSR.scala 819:37 820:23 815:30]
  wire [5:0] mstatus_lo_lo_1 = {1'h1,mstatusStruct_pie_u,mstatusStruct_ie_m,mstatusStruct_ie_h,mstatusStruct_pie_s,
    mstatusStruct_ie_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 824:27]
  wire [14:0] mstatus_lo_1 = {mstatusStruct_fs,mstatusStruct_mpp,mstatusStruct_hpp,1'h0,mstatusStruct_pie_m,
    mstatusStruct_pie_h,mstatus_lo_lo_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 824:27]
  wire [6:0] mstatus_hi_lo_1 = {mstatusStruct_tw,mstatusStruct_tvm,mstatusStruct_mxr,mstatusStruct_sum,mstatusNew_1_mprv
    ,mstatusStruct_xs}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 824:27]
  wire [63:0] _mstatus_T_9 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0
    ,mstatusStruct_tsr,mstatus_hi_lo_1,mstatus_lo_1}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 824:27]
  wire [5:0] mstatus_lo_lo_2 = {mstatusStruct_pie_s,1'h1,mstatusStruct_ie_m,mstatusStruct_ie_h,mstatusStruct_ie_s,
    mstatusStruct_pie_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 836:27]
  wire [14:0] mstatus_lo_2 = {mstatusStruct_fs,mstatusStruct_mpp,mstatusStruct_hpp,mstatusStruct_spp,mstatusStruct_pie_m
    ,mstatusStruct_pie_h,mstatus_lo_lo_2}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 836:27]
  wire [6:0] mstatus_hi_lo_2 = {mstatusStruct_tw,mstatusStruct_tvm,mstatusStruct_mxr,mstatusStruct_sum,
    mstatusStruct_mprv,mstatusStruct_xs}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 836:27]
  wire [63:0] _mstatus_T_10 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,
    mstatusStruct_pad0,mstatusStruct_tsr,mstatus_hi_lo_2,mstatus_lo_2}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 836:27]
  wire  tvalZeroWen = ~(isPageFault | isAddrMisAligned | isAccessFault) | raiseIntr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 840:73]
  wire [1:0] _GEN_60 = delegS ? priviledgeMode : {{1'd0}, mstatusStruct_spp}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19 848:22 843:30]
  wire  mstatusNew_3_pie_s = delegS ? mstatusStruct_ie_s : mstatusStruct_pie_s; // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19 849:24 843:30]
  wire  mstatusNew_3_ie_s = delegS ? 1'h0 : mstatusStruct_ie_s; // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19 850:23 843:30]
  wire [1:0] mstatusNew_3_mpp = delegS ? mstatusStruct_mpp : priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19 843:30 860:22]
  wire  mstatusNew_3_pie_m = delegS ? mstatusStruct_pie_m : mstatusStruct_ie_m; // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19 843:30 861:24]
  wire  mstatusNew_3_ie_m = delegS & mstatusStruct_ie_m; // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19 843:30 862:23]
  wire [5:0] mstatus_lo_lo_3 = {mstatusNew_3_pie_s,mstatusStruct_pie_u,mstatusNew_3_ie_m,mstatusStruct_ie_h,
    mstatusNew_3_ie_s,mstatusStruct_ie_u}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 876:27]
  wire  mstatusNew_3_spp = _GEN_60[0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 843:30]
  wire [14:0] mstatus_lo_3 = {mstatusStruct_fs,mstatusNew_3_mpp,mstatusStruct_hpp,mstatusNew_3_spp,mstatusNew_3_pie_m,
    mstatusStruct_pie_h,mstatus_lo_lo_3}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 876:27]
  wire [63:0] _mstatus_T_11 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,
    mstatusStruct_pad0,mstatusStruct_tsr,mstatus_hi_lo_2,mstatus_lo_3}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 876:27]
  wire  perfCntCondDisable_0 = wen & _T_79 & ~isIllegalMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1010:42]
  wire  _WIRE = 1'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1001:{33,33}]
  wire [63:0] _perfCnts_0_T_5 = perfCnts_0 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 986:105]
  wire  perfCntCondDisable_2 = wen & _T_81 & ~isIllegalMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1010:42]
  wire [63:0] _perfCnts_2_T_5 = perfCnts_2 + 64'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 986:105]
  wire [63:0] _perfCnts_2_T_7 = perfCnts_2 + 64'h2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 994:86]
  wire [3:0] _T_198 = raiseIntr & io_instrValid ? intrNO : 4'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1087:43]
  wire [3:0] _T_200 = raiseException & io_instrValid ? exceptionNO : 4'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1088:43]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [1:0] priviledgeMode_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:31]
  wire [1:0] priviledgeMode_t = priviledgeMode ^ priviledgeMode_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:31]
  wire  toggle_3927_clock;
  wire  toggle_3927_reset;
  wire [1:0] toggle_3927_valid;
  reg [1:0] toggle_3927_valid_reg;
  reg [63:0] mtvec_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
  wire [63:0] mtvec_t = mtvec ^ mtvec_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
  wire  toggle_3929_clock;
  wire  toggle_3929_reset;
  wire [63:0] toggle_3929_valid;
  reg [63:0] toggle_3929_valid_reg;
  reg [63:0] mcounteren_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
  wire [63:0] mcounteren_t = mcounteren ^ mcounteren_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
  wire  toggle_3993_clock;
  wire  toggle_3993_reset;
  wire [63:0] toggle_3993_valid;
  reg [63:0] toggle_3993_valid_reg;
  reg [63:0] mcause_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
  wire [63:0] mcause_t = mcause ^ mcause_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
  wire  toggle_4057_clock;
  wire  toggle_4057_reset;
  wire [63:0] toggle_4057_valid;
  reg [63:0] toggle_4057_valid_reg;
  reg [63:0] mtval_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
  wire [63:0] mtval_t = mtval ^ mtval_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
  wire  toggle_4121_clock;
  wire  toggle_4121_reset;
  wire [63:0] toggle_4121_valid;
  reg [63:0] toggle_4121_valid_reg;
  reg [63:0] mepc_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
  wire [63:0] mepc_t = mepc ^ mepc_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
  wire  toggle_4185_clock;
  wire  toggle_4185_reset;
  wire [63:0] toggle_4185_valid;
  reg [63:0] toggle_4185_valid_reg;
  reg [63:0] mie_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
  wire [63:0] mie_t = mie ^ mie_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
  wire  toggle_4249_clock;
  wire  toggle_4249_reset;
  wire [63:0] toggle_4249_valid;
  reg [63:0] toggle_4249_valid_reg;
  reg [63:0] mipReg_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
  wire [63:0] mipReg_t = mipReg ^ mipReg_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
  wire  toggle_4313_clock;
  wire  toggle_4313_reset;
  wire [63:0] toggle_4313_valid;
  reg [63:0] toggle_4313_valid_reg;
  reg [63:0] mstatus_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
  wire [63:0] mstatus_t = mstatus ^ mstatus_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
  wire  toggle_4377_clock;
  wire  toggle_4377_reset;
  wire [63:0] toggle_4377_valid;
  reg [63:0] toggle_4377_valid_reg;
  reg [63:0] medeleg_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
  wire [63:0] medeleg_t = medeleg ^ medeleg_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
  wire  toggle_4441_clock;
  wire  toggle_4441_reset;
  wire [63:0] toggle_4441_valid;
  reg [63:0] toggle_4441_valid_reg;
  reg [63:0] mideleg_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
  wire [63:0] mideleg_t = mideleg ^ mideleg_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
  wire  toggle_4505_clock;
  wire  toggle_4505_reset;
  wire [63:0] toggle_4505_valid;
  reg [63:0] toggle_4505_valid_reg;
  reg [63:0] mscratch_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
  wire [63:0] mscratch_t = mscratch ^ mscratch_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
  wire  toggle_4569_clock;
  wire  toggle_4569_reset;
  wire [63:0] toggle_4569_valid;
  reg [63:0] toggle_4569_valid_reg;
  reg [63:0] stvec_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
  wire [63:0] stvec_t = stvec ^ stvec_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
  wire  toggle_4633_clock;
  wire  toggle_4633_reset;
  wire [63:0] toggle_4633_valid;
  reg [63:0] toggle_4633_valid_reg;
  reg [63:0] satp_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
  wire [63:0] satp_t = satp ^ satp_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
  wire  toggle_4697_clock;
  wire  toggle_4697_reset;
  wire [63:0] toggle_4697_valid;
  reg [63:0] toggle_4697_valid_reg;
  reg [63:0] sepc_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
  wire [63:0] sepc_t = sepc ^ sepc_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
  wire  toggle_4761_clock;
  wire  toggle_4761_reset;
  wire [63:0] toggle_4761_valid;
  reg [63:0] toggle_4761_valid_reg;
  reg [63:0] scause_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
  wire [63:0] scause_t = scause ^ scause_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
  wire  toggle_4825_clock;
  wire  toggle_4825_reset;
  wire [63:0] toggle_4825_valid;
  reg [63:0] toggle_4825_valid_reg;
  reg [63:0] stval_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
  wire [63:0] stval_t = stval ^ stval_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
  wire  toggle_4889_clock;
  wire  toggle_4889_reset;
  wire [63:0] toggle_4889_valid;
  reg [63:0] toggle_4889_valid_reg;
  reg [63:0] sscratch_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
  wire [63:0] sscratch_t = sscratch ^ sscratch_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
  wire  toggle_4953_clock;
  wire  toggle_4953_reset;
  wire [63:0] toggle_4953_valid;
  reg [63:0] toggle_4953_valid_reg;
  reg [63:0] scounteren_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
  wire [63:0] scounteren_t = scounteren ^ scounteren_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
  wire  toggle_5017_clock;
  wire  toggle_5017_reset;
  wire [63:0] toggle_5017_valid;
  reg [63:0] toggle_5017_valid_reg;
  reg  lr_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 407:19]
  wire  lr_t = lr ^ lr_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 407:19]
  wire  toggle_5081_clock;
  wire  toggle_5081_reset;
  wire  toggle_5081_valid;
  reg  toggle_5081_valid_reg;
  reg [63:0] lrAddr_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
  wire [63:0] lrAddr_t = lrAddr ^ lrAddr_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
  wire  toggle_5082_clock;
  wire  toggle_5082_reset;
  wire [63:0] toggle_5082_valid;
  reg [63:0] toggle_5082_valid_reg;
  reg [63:0] perfCnts_0_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
  wire [63:0] perfCnts_0_t = perfCnts_0 ^ perfCnts_0_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
  wire  toggle_5146_clock;
  wire  toggle_5146_reset;
  wire [63:0] toggle_5146_valid;
  reg [63:0] toggle_5146_valid_reg;
  reg [63:0] perfCnts_1_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
  wire [63:0] perfCnts_1_t = perfCnts_1 ^ perfCnts_1_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
  wire  toggle_5210_clock;
  wire  toggle_5210_reset;
  wire [63:0] toggle_5210_valid;
  reg [63:0] toggle_5210_valid_reg;
  reg [63:0] perfCnts_2_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
  wire [63:0] perfCnts_2_t = perfCnts_2 ^ perfCnts_2_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
  wire  toggle_5274_clock;
  wire  toggle_5274_reset;
  wire [63:0] toggle_5274_valid;
  reg [63:0] toggle_5274_valid_reg;
  reg [63:0] redirectTargetReg_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
  wire [63:0] redirectTargetReg_t = redirectTargetReg ^ redirectTargetReg_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
  wire  toggle_5338_clock;
  wire  toggle_5338_reset;
  wire [63:0] toggle_5338_valid;
  reg [63:0] toggle_5338_valid_reg;
  reg  hasIllegalXRET_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 738:31]
  wire  hasIllegalXRET_t = hasIllegalXRET ^ hasIllegalXRET_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 738:31]
  wire  toggle_5402_clock;
  wire  toggle_5402_reset;
  wire  toggle_5402_valid;
  reg  toggle_5402_valid_reg;
  reg  isIllegalXRET_REG_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 739:30]
  wire  isIllegalXRET_REG_t = isIllegalXRET_REG ^ isIllegalXRET_REG_p; // @[src/main/scala/nutcore/backend/fu/CSR.scala 739:30]
  wire  toggle_5403_clock;
  wire  toggle_5403_reset;
  wire  toggle_5403_valid;
  reg  toggle_5403_valid_reg;
  CSRDiffWrapper CSRDiffWrapper ( // @[src/main/scala/nutcore/backend/fu/CSR.scala 1062:29]
    .clock(CSRDiffWrapper_clock),
    .reset(CSRDiffWrapper_reset),
    .io_csrState_privilegeMode(CSRDiffWrapper_io_csrState_privilegeMode),
    .io_csrState_mstatus(CSRDiffWrapper_io_csrState_mstatus),
    .io_csrState_sstatus(CSRDiffWrapper_io_csrState_sstatus),
    .io_csrState_mepc(CSRDiffWrapper_io_csrState_mepc),
    .io_csrState_sepc(CSRDiffWrapper_io_csrState_sepc),
    .io_csrState_mtval(CSRDiffWrapper_io_csrState_mtval),
    .io_csrState_stval(CSRDiffWrapper_io_csrState_stval),
    .io_csrState_mtvec(CSRDiffWrapper_io_csrState_mtvec),
    .io_csrState_stvec(CSRDiffWrapper_io_csrState_stvec),
    .io_csrState_mcause(CSRDiffWrapper_io_csrState_mcause),
    .io_csrState_scause(CSRDiffWrapper_io_csrState_scause),
    .io_csrState_satp(CSRDiffWrapper_io_csrState_satp),
    .io_csrState_mip(CSRDiffWrapper_io_csrState_mip),
    .io_csrState_mie(CSRDiffWrapper_io_csrState_mie),
    .io_csrState_mscratch(CSRDiffWrapper_io_csrState_mscratch),
    .io_csrState_sscratch(CSRDiffWrapper_io_csrState_sscratch),
    .io_csrState_mideleg(CSRDiffWrapper_io_csrState_mideleg),
    .io_csrState_medeleg(CSRDiffWrapper_io_csrState_medeleg),
    .io_archEvent_valid(CSRDiffWrapper_io_archEvent_valid),
    .io_archEvent_interrupt(CSRDiffWrapper_io_archEvent_interrupt),
    .io_archEvent_exception(CSRDiffWrapper_io_archEvent_exception),
    .io_archEvent_exceptionPC(CSRDiffWrapper_io_archEvent_exceptionPC),
    .io_archEvent_exceptionInst(CSRDiffWrapper_io_archEvent_exceptionInst)
  );
  GEN_w2_toggle #(.COVER_INDEX(3927)) toggle_3927 (
    .clock(toggle_3927_clock),
    .reset(toggle_3927_reset),
    .valid(toggle_3927_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(3929)) toggle_3929 (
    .clock(toggle_3929_clock),
    .reset(toggle_3929_reset),
    .valid(toggle_3929_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(3993)) toggle_3993 (
    .clock(toggle_3993_clock),
    .reset(toggle_3993_reset),
    .valid(toggle_3993_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(4057)) toggle_4057 (
    .clock(toggle_4057_clock),
    .reset(toggle_4057_reset),
    .valid(toggle_4057_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(4121)) toggle_4121 (
    .clock(toggle_4121_clock),
    .reset(toggle_4121_reset),
    .valid(toggle_4121_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(4185)) toggle_4185 (
    .clock(toggle_4185_clock),
    .reset(toggle_4185_reset),
    .valid(toggle_4185_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(4249)) toggle_4249 (
    .clock(toggle_4249_clock),
    .reset(toggle_4249_reset),
    .valid(toggle_4249_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(4313)) toggle_4313 (
    .clock(toggle_4313_clock),
    .reset(toggle_4313_reset),
    .valid(toggle_4313_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(4377)) toggle_4377 (
    .clock(toggle_4377_clock),
    .reset(toggle_4377_reset),
    .valid(toggle_4377_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(4441)) toggle_4441 (
    .clock(toggle_4441_clock),
    .reset(toggle_4441_reset),
    .valid(toggle_4441_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(4505)) toggle_4505 (
    .clock(toggle_4505_clock),
    .reset(toggle_4505_reset),
    .valid(toggle_4505_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(4569)) toggle_4569 (
    .clock(toggle_4569_clock),
    .reset(toggle_4569_reset),
    .valid(toggle_4569_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(4633)) toggle_4633 (
    .clock(toggle_4633_clock),
    .reset(toggle_4633_reset),
    .valid(toggle_4633_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(4697)) toggle_4697 (
    .clock(toggle_4697_clock),
    .reset(toggle_4697_reset),
    .valid(toggle_4697_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(4761)) toggle_4761 (
    .clock(toggle_4761_clock),
    .reset(toggle_4761_reset),
    .valid(toggle_4761_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(4825)) toggle_4825 (
    .clock(toggle_4825_clock),
    .reset(toggle_4825_reset),
    .valid(toggle_4825_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(4889)) toggle_4889 (
    .clock(toggle_4889_clock),
    .reset(toggle_4889_reset),
    .valid(toggle_4889_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(4953)) toggle_4953 (
    .clock(toggle_4953_clock),
    .reset(toggle_4953_reset),
    .valid(toggle_4953_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(5017)) toggle_5017 (
    .clock(toggle_5017_clock),
    .reset(toggle_5017_reset),
    .valid(toggle_5017_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(5081)) toggle_5081 (
    .clock(toggle_5081_clock),
    .reset(toggle_5081_reset),
    .valid(toggle_5081_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(5082)) toggle_5082 (
    .clock(toggle_5082_clock),
    .reset(toggle_5082_reset),
    .valid(toggle_5082_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(5146)) toggle_5146 (
    .clock(toggle_5146_clock),
    .reset(toggle_5146_reset),
    .valid(toggle_5146_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(5210)) toggle_5210 (
    .clock(toggle_5210_clock),
    .reset(toggle_5210_reset),
    .valid(toggle_5210_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(5274)) toggle_5274 (
    .clock(toggle_5274_clock),
    .reset(toggle_5274_reset),
    .valid(toggle_5274_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(5338)) toggle_5338 (
    .clock(toggle_5338_clock),
    .reset(toggle_5338_reset),
    .valid(toggle_5338_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(5402)) toggle_5402 (
    .clock(toggle_5402_clock),
    .reset(toggle_5402_reset),
    .valid(toggle_5402_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(5403)) toggle_5403 (
    .clock(toggle_5403_clock),
    .reset(toggle_5403_reset),
    .valid(toggle_5403_valid)
  );
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 880:16]
  assign io_out_bits = _rdata_T_113 | _rdata_T_86; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_redirect_target = redirectTarget[38:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 729:22]
  assign io_redirect_valid = io_in_valid & _isEbreak_T_1 | raiseExceptionIntr | resetSatp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 727:80]
  assign io_xretIsIllegal_valid = hasIllegalXRET; // @[src/main/scala/nutcore/backend/fu/CSR.scala 745:26]
  assign io_xretIsIllegal_bits = redirectTargetReg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 746:25]
  assign io_imemMMU_priviledgeMode = priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 603:29]
  assign io_dmemMMU_priviledgeMode = mstatusStruct_mprv ? mstatusStruct_mpp : priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 604:35]
  assign io_dmemMMU_status_sum = mstatus[18]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  assign io_dmemMMU_status_mxr = mstatus[19]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 318:39]
  assign io_wenFix = |raiseExceptionVec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 710:42]
  assign io_isPerfRead = io_out_valid & addr >= 12'hb00 & addr < 12'hb03; // @[src/main/scala/nutcore/backend/fu/CSR.scala 554:52]
  assign io_isExit = _io_isExit_T_10 & io_rfWenReal & rdata != 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 556:55]
  assign io_vmEnable = satpStruct_mode == 4'h8 & priviledgeMode < 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 251:20]
  assign io_sfence_vma_invalid = priviledgeMode == 2'h0 | tvm; // @[src/main/scala/nutcore/backend/fu/CSR.scala 542:53]
  assign io_wfi_invalid = priviledgeMode != 2'h3 & mstatusStruct_tw; // @[src/main/scala/nutcore/backend/fu/CSR.scala 546:46]
  assign lr_0 = lr;
  assign lrAddr_0 = lrAddr;
  assign satp_0 = satp;
  assign intrVecIDU_0 = intrVecIDU;
  assign CSRDiffWrapper_clock = clock;
  assign CSRDiffWrapper_reset = reset;
  assign CSRDiffWrapper_io_csrState_privilegeMode = {{62'd0}, priviledgeMode}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1066:28]
  assign CSRDiffWrapper_io_csrState_mstatus = mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1067:22]
  assign CSRDiffWrapper_io_csrState_sstatus = mstatus & 64'h80000003000d8122; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1068:33]
  assign CSRDiffWrapper_io_csrState_mepc = mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1069:19]
  assign CSRDiffWrapper_io_csrState_sepc = sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1070:19]
  assign CSRDiffWrapper_io_csrState_mtval = mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1071:19]
  assign CSRDiffWrapper_io_csrState_stval = stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1072:19]
  assign CSRDiffWrapper_io_csrState_mtvec = mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1073:20]
  assign CSRDiffWrapper_io_csrState_stvec = stvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1074:20]
  assign CSRDiffWrapper_io_csrState_mcause = mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1075:21]
  assign CSRDiffWrapper_io_csrState_scause = scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1076:21]
  assign CSRDiffWrapper_io_csrState_satp = satp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1077:19]
  assign CSRDiffWrapper_io_csrState_mip = mipReg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1078:18]
  assign CSRDiffWrapper_io_csrState_mie = mie; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1079:18]
  assign CSRDiffWrapper_io_csrState_mscratch = mscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1080:23]
  assign CSRDiffWrapper_io_csrState_sscratch = sscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1081:23]
  assign CSRDiffWrapper_io_csrState_mideleg = mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1082:22]
  assign CSRDiffWrapper_io_csrState_medeleg = medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1083:22]
  assign CSRDiffWrapper_io_archEvent_valid = (raiseException | raiseIntr) & io_instrValid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 717:58]
  assign CSRDiffWrapper_io_archEvent_interrupt = {{28'd0}, _T_198}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1087:37]
  assign CSRDiffWrapper_io_archEvent_exception = {{28'd0}, _T_200}; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1088:37]
  assign CSRDiffWrapper_io_archEvent_exceptionPC = io_illegalJump_valid ? io_illegalJump_bits : _imemExceptionAddr_T_11; // @[src/main/scala/nutcore/backend/fu/CSR.scala 648:23]
  assign CSRDiffWrapper_io_archEvent_exceptionInst = io_cfIn_instr[31:0]; // @[src/main/scala/nutcore/backend/fu/CSR.scala 1090:37]
  assign toggle_3927_clock = clock;
  assign toggle_3927_reset = reset;
  assign toggle_3927_valid = priviledgeMode ^ toggle_3927_valid_reg;
  assign toggle_3929_clock = clock;
  assign toggle_3929_reset = reset;
  assign toggle_3929_valid = mtvec ^ toggle_3929_valid_reg;
  assign toggle_3993_clock = clock;
  assign toggle_3993_reset = reset;
  assign toggle_3993_valid = mcounteren ^ toggle_3993_valid_reg;
  assign toggle_4057_clock = clock;
  assign toggle_4057_reset = reset;
  assign toggle_4057_valid = mcause ^ toggle_4057_valid_reg;
  assign toggle_4121_clock = clock;
  assign toggle_4121_reset = reset;
  assign toggle_4121_valid = mtval ^ toggle_4121_valid_reg;
  assign toggle_4185_clock = clock;
  assign toggle_4185_reset = reset;
  assign toggle_4185_valid = mepc ^ toggle_4185_valid_reg;
  assign toggle_4249_clock = clock;
  assign toggle_4249_reset = reset;
  assign toggle_4249_valid = mie ^ toggle_4249_valid_reg;
  assign toggle_4313_clock = clock;
  assign toggle_4313_reset = reset;
  assign toggle_4313_valid = mipReg ^ toggle_4313_valid_reg;
  assign toggle_4377_clock = clock;
  assign toggle_4377_reset = reset;
  assign toggle_4377_valid = mstatus ^ toggle_4377_valid_reg;
  assign toggle_4441_clock = clock;
  assign toggle_4441_reset = reset;
  assign toggle_4441_valid = medeleg ^ toggle_4441_valid_reg;
  assign toggle_4505_clock = clock;
  assign toggle_4505_reset = reset;
  assign toggle_4505_valid = mideleg ^ toggle_4505_valid_reg;
  assign toggle_4569_clock = clock;
  assign toggle_4569_reset = reset;
  assign toggle_4569_valid = mscratch ^ toggle_4569_valid_reg;
  assign toggle_4633_clock = clock;
  assign toggle_4633_reset = reset;
  assign toggle_4633_valid = stvec ^ toggle_4633_valid_reg;
  assign toggle_4697_clock = clock;
  assign toggle_4697_reset = reset;
  assign toggle_4697_valid = satp ^ toggle_4697_valid_reg;
  assign toggle_4761_clock = clock;
  assign toggle_4761_reset = reset;
  assign toggle_4761_valid = sepc ^ toggle_4761_valid_reg;
  assign toggle_4825_clock = clock;
  assign toggle_4825_reset = reset;
  assign toggle_4825_valid = scause ^ toggle_4825_valid_reg;
  assign toggle_4889_clock = clock;
  assign toggle_4889_reset = reset;
  assign toggle_4889_valid = stval ^ toggle_4889_valid_reg;
  assign toggle_4953_clock = clock;
  assign toggle_4953_reset = reset;
  assign toggle_4953_valid = sscratch ^ toggle_4953_valid_reg;
  assign toggle_5017_clock = clock;
  assign toggle_5017_reset = reset;
  assign toggle_5017_valid = scounteren ^ toggle_5017_valid_reg;
  assign toggle_5081_clock = clock;
  assign toggle_5081_reset = reset;
  assign toggle_5081_valid = lr ^ toggle_5081_valid_reg;
  assign toggle_5082_clock = clock;
  assign toggle_5082_reset = reset;
  assign toggle_5082_valid = lrAddr ^ toggle_5082_valid_reg;
  assign toggle_5146_clock = clock;
  assign toggle_5146_reset = reset;
  assign toggle_5146_valid = perfCnts_0 ^ toggle_5146_valid_reg;
  assign toggle_5210_clock = clock;
  assign toggle_5210_reset = reset;
  assign toggle_5210_valid = perfCnts_1 ^ toggle_5210_valid_reg;
  assign toggle_5274_clock = clock;
  assign toggle_5274_reset = reset;
  assign toggle_5274_valid = perfCnts_2 ^ toggle_5274_valid_reg;
  assign toggle_5338_clock = clock;
  assign toggle_5338_reset = reset;
  assign toggle_5338_valid = redirectTargetReg ^ toggle_5338_valid_reg;
  assign toggle_5402_clock = clock;
  assign toggle_5402_reset = reset;
  assign toggle_5402_valid = hasIllegalXRET ^ toggle_5402_valid_reg;
  assign toggle_5403_clock = clock;
  assign toggle_5403_reset = reset;
  assign toggle_5403_valid = isIllegalXRET_REG ^ toggle_5403_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:31]
      priviledgeMode <= 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:31]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19]
        priviledgeMode <= 2'h1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 851:22]
      end else begin
        priviledgeMode <= 2'h3; // @[src/main/scala/nutcore/backend/fu/CSR.scala 863:22]
      end
    end else if (io_in_valid & isUret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 829:26]
      priviledgeMode <= 2'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 834:20]
    end else if (_illegalSret_T & ~illegalSret & ~illegalSModeSret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 813:63]
      priviledgeMode <= _priviledgeMode_T; // @[src/main/scala/nutcore/backend/fu/CSR.scala 818:20]
    end else begin
      priviledgeMode <= _GEN_44;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
      mtvec <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end else if (canWriteCSR & addr == 12'h305) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mtvec <= _mtvec_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
      mcounteren <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end else if (canWriteCSR & addr == 12'h306) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mcounteren <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
      mcause <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19]
        mcause <= _GEN_14;
      end else begin
        mcause <= causeNO; // @[src/main/scala/nutcore/backend/fu/CSR.scala 858:14]
      end
    end else begin
      mcause <= _GEN_14;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
      mtval <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19]
        mtval <= _GEN_42;
      end else if (tvalZeroWen) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 864:26]
        mtval <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 865:15]
      end else begin
        mtval <= _GEN_42;
      end
    end else begin
      mtval <= _GEN_42;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
      mepc <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19]
        mepc <= _GEN_21;
      end else if (io_illegalJump_valid) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 648:23]
        mepc <= io_illegalJump_bits;
      end else begin
        mepc <= _imemExceptionAddr_T_11;
      end
    end else begin
      mepc <= _GEN_21;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
      mie <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end else if (canWriteCSR & addr == 12'h304) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mie <= _mie_T_7; // @[src/main/scala/utils/RegMap.scala 50:76]
    end else if (canWriteCSR & addr == 12'h104) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mie <= _mie_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
      mipReg <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end else if (_canWriteCSR_T_1 & _io_isExit_T_1) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mipReg <= _mipReg_T_7; // @[src/main/scala/utils/RegMap.scala 50:76]
    end else if (_canWriteCSR_T_1 & _io_isExit_T) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mipReg <= _mipReg_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
      mstatus <= 64'ha00001800; // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:29]
      mstatus <= _mstatus_T_11; // @[src/main/scala/nutcore/backend/fu/CSR.scala 876:13]
    end else if (io_in_valid & isUret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 829:26]
      mstatus <= _mstatus_T_10; // @[src/main/scala/nutcore/backend/fu/CSR.scala 836:13]
    end else if (_illegalSret_T & ~illegalSret & ~illegalSModeSret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 813:63]
      mstatus <= _mstatus_T_9; // @[src/main/scala/nutcore/backend/fu/CSR.scala 824:13]
    end else begin
      mstatus <= _GEN_45;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
      medeleg <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end else if (canWriteCSR & addr == 12'h302) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      medeleg <= _medeleg_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
      mideleg <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end else if (canWriteCSR & addr == 12'h303) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mideleg <= _mideleg_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
      mscratch <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end else if (canWriteCSR & addr == 12'h340) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      mscratch <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
      stvec <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end else if (canWriteCSR & addr == 12'h105) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      stvec <= _stvec_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
      satp <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end else if (canWriteCSR & _isIllegalTVM_T_1) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      satp <= _satp_T_3; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
      sepc <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19]
        if (io_illegalJump_valid) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 648:23]
          sepc <= io_illegalJump_bits;
        end else begin
          sepc <= _imemExceptionAddr_T_11;
        end
      end else begin
        sepc <= _GEN_13;
      end
    end else begin
      sepc <= _GEN_13;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
      scause <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19]
        scause <= causeNO; // @[src/main/scala/nutcore/backend/fu/CSR.scala 846:14]
      end else begin
        scause <= _GEN_10;
      end
    end else begin
      scause <= _GEN_10;
    end
    if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 841:29]
      if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 845:19]
        if (tvalZeroWen) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 852:26]
          stval <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 853:15]
        end else begin
          stval <= _GEN_41;
        end
      end else begin
        stval <= _GEN_41;
      end
    end else begin
      stval <= _GEN_41;
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
      sscratch <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end else if (canWriteCSR & addr == 12'h140) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      sscratch <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
      scounteren <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end else if (canWriteCSR & addr == 12'h106) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      scounteren <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 407:19]
      lr <= 1'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 407:19]
    end else if (_illegalSret_T & ~illegalSret & ~illegalSModeSret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 813:63]
      lr <= 1'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 825:8]
    end else if (_illegalMret_T & ~illegalMret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 797:42]
      lr <= 1'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 809:8]
    end else if (set_lr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 415:14]
      lr <= set_lr_val; // @[src/main/scala/nutcore/backend/fu/CSR.scala 416:8]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
      lrAddr <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end else if (set_lr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 415:14]
      lrAddr <= set_lr_addr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 417:12]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
      perfCnts_0 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end else if (~perfCntCondDisable_0) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 986:96]
      perfCnts_0 <= _perfCnts_0_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 986:100]
    end else if (canWriteCSR & addr == 12'hb00) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_0 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
      perfCnts_1 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end else if (canWriteCSR & addr == 12'hb01) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_1 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
      perfCnts_2 <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end else if (perfCntCondMultiCommit) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 994:35]
      perfCnts_2 <= _perfCnts_2_T_7; // @[src/main/scala/nutcore/backend/fu/CSR.scala 994:60]
    end else if (perfCntCondMinstret & ~perfCntCondDisable_2) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 986:96]
      perfCnts_2 <= _perfCnts_2_T_5; // @[src/main/scala/nutcore/backend/fu/CSR.scala 986:100]
    end else if (canWriteCSR & addr == 12'hb02) begin // @[src/main/scala/utils/RegMap.scala 50:72]
      perfCnts_2 <= wdata; // @[src/main/scala/utils/RegMap.scala 50:76]
    end
    if (io_redirect_valid) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
      if (resetSatp) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 720:27]
        redirectTargetReg <= _redirectTarget_T_3;
      end else if (raiseExceptionIntr) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 722:8]
        if (delegS) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 766:20]
          redirectTargetReg <= stvec;
        end else begin
          redirectTargetReg <= mtvec;
        end
      end else if (io_in_valid & isUret) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 829:26]
        redirectTargetReg <= 64'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 837:15]
      end else begin
        redirectTargetReg <= _GEN_52;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/fu/CSR.scala 738:31]
      hasIllegalXRET <= 1'h0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 738:31]
    end else begin
      hasIllegalXRET <= _GEN_28;
    end
    isIllegalXRET_REG <= io_redirect_valid; // @[src/main/scala/nutcore/backend/fu/CSR.scala 739:30]
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    priviledgeMode_p <= priviledgeMode; // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:31]
    toggle_3927_valid_reg <= priviledgeMode;
    mtvec_p <= mtvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    toggle_3929_valid_reg <= mtvec;
    mcounteren_p <= mcounteren; // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    toggle_3993_valid_reg <= mcounteren;
    mcause_p <= mcause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    toggle_4057_valid_reg <= mcause;
    mtval_p <= mtval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    toggle_4121_valid_reg <= mtval;
    mepc_p <= mepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    toggle_4185_valid_reg <= mepc;
    mie_p <= mie; // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    toggle_4249_valid_reg <= mie;
    mipReg_p <= mipReg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    toggle_4313_valid_reg <= mipReg;
    mstatus_p <= mstatus; // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    toggle_4377_valid_reg <= mstatus;
    medeleg_p <= medeleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    toggle_4441_valid_reg <= medeleg;
    mideleg_p <= mideleg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    toggle_4505_valid_reg <= mideleg;
    mscratch_p <= mscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    toggle_4569_valid_reg <= mscratch;
    stvec_p <= stvec; // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    toggle_4633_valid_reg <= stvec;
    satp_p <= satp; // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    toggle_4697_valid_reg <= satp;
    sepc_p <= sepc; // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    toggle_4761_valid_reg <= sepc;
    scause_p <= scause; // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    toggle_4825_valid_reg <= scause;
    stval_p <= stval; // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    toggle_4889_valid_reg <= stval;
    sscratch_p <= sscratch; // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    toggle_4953_valid_reg <= sscratch;
    scounteren_p <= scounteren; // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    toggle_5017_valid_reg <= scounteren;
    lr_p <= lr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 407:19]
    toggle_5081_valid_reg <= lr;
    lrAddr_p <= lrAddr; // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    toggle_5082_valid_reg <= lrAddr;
    perfCnts_0_p <= perfCnts_0; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    toggle_5146_valid_reg <= perfCnts_0;
    perfCnts_1_p <= perfCnts_1; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    toggle_5210_valid_reg <= perfCnts_1;
    perfCnts_2_p <= perfCnts_2; // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    toggle_5274_valid_reg <= perfCnts_2;
    redirectTargetReg_p <= redirectTargetReg; // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    toggle_5338_valid_reg <= redirectTargetReg;
    hasIllegalXRET_p <= hasIllegalXRET; // @[src/main/scala/nutcore/backend/fu/CSR.scala 738:31]
    toggle_5402_valid_reg <= hasIllegalXRET;
    isIllegalXRET_REG_p <= isIllegalXRET_REG; // @[src/main/scala/nutcore/backend/fu/CSR.scala 739:30]
    toggle_5403_valid_reg <= isIllegalXRET_REG;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  priviledgeMode = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  mtvec = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mcounteren = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mcause = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mtval = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mepc = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mie = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  mipReg = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  mstatus = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  medeleg = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  mideleg = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  mscratch = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  stvec = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  satp = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  sepc = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  scause = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  stval = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  sscratch = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  scounteren = _RAND_18[63:0];
  _RAND_19 = {1{`RANDOM}};
  lr = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  lrAddr = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  perfCnts_0 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  perfCnts_1 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  perfCnts_2 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  redirectTargetReg = _RAND_24[63:0];
  _RAND_25 = {1{`RANDOM}};
  hasIllegalXRET = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  isIllegalXRET_REG = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  priviledgeMode_p = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  toggle_3927_valid_reg = _RAND_28[1:0];
  _RAND_29 = {2{`RANDOM}};
  mtvec_p = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  toggle_3929_valid_reg = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  mcounteren_p = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  toggle_3993_valid_reg = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  mcause_p = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  toggle_4057_valid_reg = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  mtval_p = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  toggle_4121_valid_reg = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  mepc_p = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  toggle_4185_valid_reg = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  mie_p = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  toggle_4249_valid_reg = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  mipReg_p = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  toggle_4313_valid_reg = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  mstatus_p = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  toggle_4377_valid_reg = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  medeleg_p = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  toggle_4441_valid_reg = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  mideleg_p = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  toggle_4505_valid_reg = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  mscratch_p = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  toggle_4569_valid_reg = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  stvec_p = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  toggle_4633_valid_reg = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  satp_p = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  toggle_4697_valid_reg = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  sepc_p = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  toggle_4761_valid_reg = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  scause_p = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  toggle_4825_valid_reg = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  stval_p = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  toggle_4889_valid_reg = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  sscratch_p = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  toggle_4953_valid_reg = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  scounteren_p = _RAND_63[63:0];
  _RAND_64 = {2{`RANDOM}};
  toggle_5017_valid_reg = _RAND_64[63:0];
  _RAND_65 = {1{`RANDOM}};
  lr_p = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  toggle_5081_valid_reg = _RAND_66[0:0];
  _RAND_67 = {2{`RANDOM}};
  lrAddr_p = _RAND_67[63:0];
  _RAND_68 = {2{`RANDOM}};
  toggle_5082_valid_reg = _RAND_68[63:0];
  _RAND_69 = {2{`RANDOM}};
  perfCnts_0_p = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  toggle_5146_valid_reg = _RAND_70[63:0];
  _RAND_71 = {2{`RANDOM}};
  perfCnts_1_p = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  toggle_5210_valid_reg = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  perfCnts_2_p = _RAND_73[63:0];
  _RAND_74 = {2{`RANDOM}};
  toggle_5274_valid_reg = _RAND_74[63:0];
  _RAND_75 = {2{`RANDOM}};
  redirectTargetReg_p = _RAND_75[63:0];
  _RAND_76 = {2{`RANDOM}};
  toggle_5338_valid_reg = _RAND_76[63:0];
  _RAND_77 = {1{`RANDOM}};
  hasIllegalXRET_p = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  toggle_5402_valid_reg = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  isIllegalXRET_REG_p = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  toggle_5403_valid_reg = _RAND_80[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(priviledgeMode_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:31]
    end
    //
    if (enToggle_past) begin
      cover(priviledgeMode_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 262:31]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mtvec_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 266:22]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcounteren_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 268:27]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mcause_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 269:23]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mtval_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 270:22]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mepc_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 273:21]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mie_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 276:20]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mipReg_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 279:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(mstatus_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 297:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(medeleg_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 351:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mideleg_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 352:24]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(mscratch_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 353:25]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(stvec_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 376:22]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(satp_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 382:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(sepc_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 388:21]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(scause_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 391:23]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(stval_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 392:18]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(sscratch_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 393:25]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(scounteren_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 394:27]
    end
    //
    if (enToggle_past) begin
      cover(lr_t); // @[src/main/scala/nutcore/backend/fu/CSR.scala 407:19]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(lrAddr_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 408:23]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_0_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_1_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(perfCnts_2_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 424:47]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[0]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[1]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[2]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[3]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[4]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[5]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[6]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[7]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[8]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[9]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[10]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[11]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[12]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[13]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[14]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[15]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[16]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[17]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[18]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[19]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[20]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[21]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[22]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[23]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[24]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[25]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[26]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[27]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[28]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[29]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[30]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[31]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[32]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[33]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[34]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[35]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[36]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[37]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[38]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[39]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[40]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[41]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[42]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[43]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[44]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[45]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[46]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[47]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[48]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[49]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[50]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[51]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[52]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[53]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[54]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[55]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[56]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[57]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[58]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[59]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[60]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[61]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[62]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(redirectTargetReg_t[63]); // @[src/main/scala/nutcore/backend/fu/CSR.scala 733:36]
    end
    //
    if (enToggle_past) begin
      cover(hasIllegalXRET_t); // @[src/main/scala/nutcore/backend/fu/CSR.scala 738:31]
    end
    //
    if (enToggle_past) begin
      cover(isIllegalXRET_REG_t); // @[src/main/scala/nutcore/backend/fu/CSR.scala 739:30]
    end
  end
endmodule
module MOU(
  input         clock,
  input         reset,
  input         io_in_valid, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  input  [6:0]  io_in_bits_func, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  input  [38:0] io_cfIn_pc, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  output [38:0] io_redirect_target, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  output        io_redirect_valid, // @[src/main/scala/nutcore/backend/fu/MOU.scala 38:14]
  output        flushICache_0,
  output        flushTLB_0
);
  wire  flushICache = io_in_valid & io_in_bits_func == 7'h1; // @[src/main/scala/nutcore/backend/fu/MOU.scala 52:27]
  wire  flushTLB = io_in_valid & io_in_bits_func == 7'h2; // @[src/main/scala/nutcore/backend/fu/MOU.scala 56:24]
  assign io_redirect_target = io_cfIn_pc + 39'h4; // @[src/main/scala/nutcore/backend/fu/MOU.scala 49:36]
  assign io_redirect_valid = io_in_valid; // @[src/main/scala/nutcore/backend/fu/MOU.scala 50:21]
  assign flushICache_0 = flushICache;
  assign flushTLB_0 = flushTLB;
endmodule
module DummyDPICWrapper_3(
  input         clock,
  input         reset,
  input         io_bits_hasTrap, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_cycleCnt, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_instrCnt, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [31:0] io_bits_code, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_pc // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_hasTrap; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_cycleCnt; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_instrCnt; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_hasWFI; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [31:0] dpic_io_code; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_pc; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestTrapEvent dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_hasTrap(dpic_io_hasTrap),
    .io_cycleCnt(dpic_io_cycleCnt),
    .io_instrCnt(dpic_io_instrCnt),
    .io_hasWFI(dpic_io_hasWFI),
    .io_code(dpic_io_code),
    .io_pc(dpic_io_pc),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = 1'h1; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_hasTrap = io_bits_hasTrap; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_cycleCnt = io_bits_cycleCnt; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_instrCnt = io_bits_instrCnt; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_hasWFI = 1'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_code = io_bits_code; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_pc = io_bits_pc; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module EXUDiffWrapper(
  input         clock,
  input         reset,
  input         io_in_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 179:14]
  input  [38:0] io_in_bits_cf_pc, // @[src/main/scala/nutcore/backend/seq/EXU.scala 179:14]
  input         io_in_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/backend/seq/EXU.scala 179:14]
  input  [63:0] io_in_bits_data_src1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 179:14]
  input         io_flush, // @[src/main/scala/nutcore/backend/seq/EXU.scala 179:14]
  input         perfCntCondMinstret
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  difftest_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_hasTrap; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_cycleCnt; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_instrCnt; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [31:0] difftest_module_io_bits_code; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_pc; // @[difftest/src/main/scala/DPIC.scala 299:24]
  reg [63:0] cycleCnt; // @[src/main/scala/nutcore/backend/seq/EXU.scala 185:25]
  wire [63:0] _cycleCnt_T_1 = cycleCnt + 64'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 186:24]
  reg [63:0] instrCnt; // @[src/main/scala/nutcore/backend/seq/EXU.scala 187:25]
  wire [63:0] _instrCnt_T_1 = instrCnt + 64'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 190:26]
  wire  nutcoretrap = io_in_bits_ctrl_isNutCoreTrap & io_in_valid & ~io_flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 194:66]
  DummyDPICWrapper_3 difftest_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_clock),
    .reset(difftest_module_reset),
    .io_bits_hasTrap(difftest_module_io_bits_hasTrap),
    .io_bits_cycleCnt(difftest_module_io_bits_cycleCnt),
    .io_bits_instrCnt(difftest_module_io_bits_instrCnt),
    .io_bits_code(difftest_module_io_bits_code),
    .io_bits_pc(difftest_module_io_bits_pc)
  );
  assign difftest_module_clock = clock;
  assign difftest_module_reset = reset;
  assign difftest_module_io_bits_hasTrap = nutcoretrap; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/EXU.scala 199:21]
  assign difftest_module_io_bits_cycleCnt = cycleCnt; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/EXU.scala 202:21]
  assign difftest_module_io_bits_instrCnt = instrCnt; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/EXU.scala 203:21]
  assign difftest_module_io_bits_code = io_in_bits_data_src1[31:0]; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/EXU.scala 200:21]
  assign difftest_module_io_bits_pc = {{25'd0}, io_in_bits_cf_pc}; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/EXU.scala 201:21]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 185:25]
      cycleCnt <= 64'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 185:25]
    end else begin
      cycleCnt <= _cycleCnt_T_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 186:12]
    end
    if (reset) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 187:25]
      instrCnt <= 64'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 187:25]
    end else if (perfCntCondMinstret) begin // @[src/main/scala/nutcore/backend/seq/EXU.scala 189:22]
      instrCnt <= _instrCnt_T_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 190:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  cycleCnt = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  instrCnt = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EXU(
  input         clock,
  input         reset,
  output        io__in_ready, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [63:0] io__in_bits_cf_instr, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [38:0] io__in_bits_cf_pc, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [38:0] io__in_bits_cf_pnpc, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_intrVec_1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_intrVec_3, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_intrVec_5, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_intrVec_7, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_intrVec_9, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_intrVec_11, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [3:0]  io__in_bits_cf_brIdx, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [2:0]  io__in_bits_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [6:0]  io__in_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [4:0]  io__in_bits_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__in_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [63:0] io__in_bits_data_src1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [63:0] io__in_bits_data_src2, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [63:0] io__in_bits_data_imm, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__out_ready, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__out_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__out_bits_decode_cf_instr, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [38:0] io__out_bits_decode_cf_pc, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [38:0] io__out_bits_decode_cf_redirect_target, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__out_bits_decode_cf_redirect_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [2:0]  io__out_bits_decode_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__out_bits_decode_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [4:0]  io__out_bits_decode_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__out_bits_isMMIO, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__out_bits_commits_0, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__out_bits_commits_1, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__out_bits_commits_2, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__out_bits_commits_3, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__out_bits_isExit, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__flush, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__dmem_req_ready, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__dmem_req_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [38:0] io__dmem_req_bits_addr, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [2:0]  io__dmem_req_bits_size, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [3:0]  io__dmem_req_bits_cmd, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [7:0]  io__dmem_req_bits_wmask, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__dmem_req_bits_wdata, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__dmem_resp_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input  [63:0] io__dmem_resp_bits_rdata, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__forward_valid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__forward_wb_rfWen, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [4:0]  io__forward_wb_rfDest, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [63:0] io__forward_wb_rfData, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [2:0]  io__forward_fuType, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [1:0]  io__memMMU_imem_priviledgeMode, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output [1:0]  io__memMMU_dmem_priviledgeMode, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__memMMU_dmem_status_sum, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__memMMU_dmem_status_mxr, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__memMMU_dmem_loadPF, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__memMMU_dmem_storePF, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__memMMU_dmem_laf, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  input         io__memMMU_dmem_saf, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__sfence_vma_invalid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        io__wfi_invalid, // @[src/main/scala/nutcore/backend/seq/EXU.scala 30:14]
  output        lr,
  input         io_extra_meip_0,
  output        scInflight,
  output        REG_valid,
  output [38:0] REG_pc,
  output        REG_isMissPredict,
  output [38:0] REG_actualTarget,
  output [6:0]  REG_fuOpType,
  output [1:0]  REG_btbType,
  output        REG_isRVC,
  output        amoReq,
  output [63:0] lrAddr,
  input  [55:0] paddr,
  output [63:0] satp,
  input         _T_12_0,
  input         scIsSuccess,
  input         io_extra_mtip,
  output        flushICache,
  input         falseWire,
  input         vmEnable,
  output        flushTLB,
  output [11:0] intrVecIDU,
  input         tlbFinish,
  input         ismmio,
  input         _T_13_1,
  input         io_extra_msip,
  input         io_in_valid
);
  wire  alu_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [63:0] alu_io_in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [63:0] alu_io_in_bits_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [6:0] alu_io_in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_out_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [63:0] alu_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [63:0] alu_io_cfIn_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [38:0] alu_io_cfIn_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [38:0] alu_io_cfIn_pnpc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [3:0] alu_io_cfIn_brIdx; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [38:0] alu_io_redirect_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [63:0] alu_io_offset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_iVmEnable; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_jumpIsIllegal_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_io_jumpIsIllegal_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [63:0] alu_io_jumpIsIllegal_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_REG_0_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [38:0] alu_REG_0_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_REG_0_isMissPredict; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [38:0] alu_REG_0_actualTarget; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [6:0] alu_REG_0_fuOpType; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire [1:0] alu_REG_0_btbType; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  alu_REG_0_isRVC; // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
  wire  lsu_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__in_bits_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [6:0] lsu_io__in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__out_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__wdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [31:0] lsu_io__instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__dmem_req_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [38:0] lsu_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [2:0] lsu_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [3:0] lsu_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [7:0] lsu_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__isMMIO; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__dtlbPF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__dtlbAF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_io__vaddr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__loadAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__storeAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__loadAccessFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_io__storeAccessFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_setLr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_lr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_scInflight_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_amoReq_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_lr_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [55:0] lsu_dtlb_paddr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu__T_12_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_scIsSuccess_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_setLrVal_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_vmEnable; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_DTLBFINISH; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu_lsuMMIO_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  lsu__T_13_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire [63:0] lsu_setLrAddr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
  wire  mdu_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire  mdu_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire  mdu_io_in_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire  mdu_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire [63:0] mdu_io_in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire [63:0] mdu_io_in_bits_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire [6:0] mdu_io_in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire  mdu_io_out_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire  mdu_io_out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire [63:0] mdu_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
  wire  csr_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_in_bits_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_in_bits_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [6:0] csr_io_in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_out_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_cfIn_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [38:0] csr_io_cfIn_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_4; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_5; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_6; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_7; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_12; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_13; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_exceptionVec_15; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_intrVec_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_intrVec_3; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_intrVec_5; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_intrVec_7; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_intrVec_9; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_intrVec_11; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_cfIn_crossBoundaryFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [38:0] csr_io_redirect_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_instrValid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_illegalJump_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_illegalJump_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_dmemExceptionAddr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_xretIsIllegal_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_xretIsIllegal_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_io_xretIsIllegal_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [1:0] csr_io_imemMMU_priviledgeMode; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [1:0] csr_io_dmemMMU_priviledgeMode; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_dmemMMU_status_sum; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_dmemMMU_status_mxr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_dmemMMU_loadPF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_dmemMMU_storePF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_dmemMMU_laf; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_dmemMMU_saf; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_wenFix; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_isPerfRead; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_isExit; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_vmEnable; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_rfWenReal; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_sfence_vma_invalid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_io_wfi_invalid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_set_lr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_lr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_meip_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_lrAddr_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_satp_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_mtip_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_perfCntCondMultiCommit; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_set_lr_val; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [11:0] csr_intrVecIDU_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire [63:0] csr_set_lr_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_msip_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  csr_perfCntCondMinstret; // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
  wire  mou_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire  mou_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire  mou_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire [6:0] mou_io_in_bits_func; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire [38:0] mou_io_cfIn_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire [38:0] mou_io_redirect_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire  mou_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire  mou_flushICache_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire  mou_flushTLB_0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
  wire  diffMod_clock; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire  diffMod_reset; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire  diffMod_io_in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire [38:0] diffMod_io_in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire  diffMod_io_in_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire [63:0] diffMod_io_in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire  diffMod_io_flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire  diffMod_perfCntCondMinstret; // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
  wire  _fuValids_0_T_2 = ~io__flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 47:84]
  wire [15:0] _fuValids_0_T_4 = {2'h0,1'h0,io__in_bits_cf_exceptionVec_12,4'h0,4'h0,1'h0,io__in_bits_cf_exceptionVec_2,
    io__in_bits_cf_exceptionVec_1,1'h0}; // @[src/main/scala/nutcore/backend/seq/EXU.scala 47:125]
  wire  _csr_io_cfIn_exceptionVec_13_T = lsu_io__in_valid & lsu_io__dtlbPF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 78:62]
  wire  _csr_io_cfIn_exceptionVec_13_T_2 = io__in_bits_ctrl_fuOpType == 7'h20; // @[src/main/scala/nutcore/backend/fu/LSU.scala 57:37]
  wire  _csr_io_cfIn_exceptionVec_13_T_6 = io__in_bits_ctrl_fuOpType[5] & ~_csr_io_cfIn_exceptionVec_13_T_2 |
    io__in_bits_ctrl_fuOpType[3]; // @[src/main/scala/nutcore/backend/fu/LSU.scala 64:69]
  wire  _csr_io_cfIn_exceptionVec_13_T_7 = ~_csr_io_cfIn_exceptionVec_13_T_6; // @[src/main/scala/nutcore/backend/fu/LSU.scala 65:40]
  wire  _T = alu_io_jumpIsIllegal_ready & alu_io_jumpIsIllegal_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_1 = csr_io_xretIsIllegal_ready & csr_io_xretIsIllegal_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _GEN_0 = csr_io_vmEnable | io__in_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/seq/EXU.scala 103:28 104:48 73:15]
  wire  _GEN_1 = csr_io_vmEnable ? io__in_bits_cf_exceptionVec_1 : 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 103:28 73:15 106:50]
  wire  fuValids_1 = _T | _T_1 ? 1'h0 : io__in_bits_ctrl_fuType == 3'h1 & io__in_valid & ~io__flush & ~(|_fuValids_0_T_4
    ); // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  wire  fuValids_3 = _T | _T_1 | io__in_bits_ctrl_fuType == 3'h3 & io__in_valid & ~io__flush & ~(|_fuValids_0_T_4); // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  wire  lsuTlbPF = lsu_io__dtlbPF; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 53:12 src/main/scala/nutcore/backend/seq/EXU.scala 58:26]
  wire  _hasException_T_1 = lsuTlbPF | lsu_io__dtlbAF | lsu_io__loadAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 123:50]
  wire  _hasException_T_3 = _hasException_T_1 | lsu_io__storeAddrMisaligned | lsu_io__loadAccessFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 124:63]
  wire  hasException = _hasException_T_3 | lsu_io__storeAccessFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 125:30]
  wire [38:0] _io_out_bits_decode_cf_redirect_T_target = csr_io_redirect_valid ? csr_io_redirect_target :
    alu_io_redirect_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 137:10]
  wire  _io_out_bits_decode_cf_redirect_T_valid = csr_io_redirect_valid ? csr_io_redirect_valid : alu_io_redirect_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 137:10]
  wire  _io_out_valid_T_1 = 3'h1 == io__in_bits_ctrl_fuType ? lsu_io__out_valid : 1'h1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _io_out_valid_T_3 = 3'h2 == io__in_bits_ctrl_fuType ? mdu_io_out_valid : _io_out_valid_T_1; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _io_out_valid_T_4 = _io_out_valid_T_3 | csr_io_illegalJump_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 146:6]
  wire  _io_forward_wb_rfData_T = alu_io_out_ready & alu_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  isBru = io__in_bits_ctrl_fuOpType[4]; // @[src/main/scala/nutcore/backend/fu/ALU.scala 62:31]
  wire  _T_10 = _io_forward_wb_rfData_T & ~isBru; // @[src/main/scala/nutcore/backend/seq/EXU.scala 163:43]
  wire  _T_12 = _io_forward_wb_rfData_T & isBru; // @[src/main/scala/nutcore/backend/seq/EXU.scala 164:43]
  wire  _T_13 = lsu_io__out_ready & lsu_io__out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_14 = mdu_io_out_ready & mdu_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_15 = csr_io_out_ready & csr_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  ALU alu ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 49:19]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_in_valid(alu_io_in_valid),
    .io_in_bits_src1(alu_io_in_bits_src1),
    .io_in_bits_src2(alu_io_in_bits_src2),
    .io_in_bits_func(alu_io_in_bits_func),
    .io_out_ready(alu_io_out_ready),
    .io_out_valid(alu_io_out_valid),
    .io_out_bits(alu_io_out_bits),
    .io_cfIn_instr(alu_io_cfIn_instr),
    .io_cfIn_pc(alu_io_cfIn_pc),
    .io_cfIn_pnpc(alu_io_cfIn_pnpc),
    .io_cfIn_brIdx(alu_io_cfIn_brIdx),
    .io_redirect_target(alu_io_redirect_target),
    .io_redirect_valid(alu_io_redirect_valid),
    .io_offset(alu_io_offset),
    .io_iVmEnable(alu_io_iVmEnable),
    .io_jumpIsIllegal_ready(alu_io_jumpIsIllegal_ready),
    .io_jumpIsIllegal_valid(alu_io_jumpIsIllegal_valid),
    .io_jumpIsIllegal_bits(alu_io_jumpIsIllegal_bits),
    .REG_0_valid(alu_REG_0_valid),
    .REG_0_pc(alu_REG_0_pc),
    .REG_0_isMissPredict(alu_REG_0_isMissPredict),
    .REG_0_actualTarget(alu_REG_0_actualTarget),
    .REG_0_fuOpType(alu_REG_0_fuOpType),
    .REG_0_btbType(alu_REG_0_btbType),
    .REG_0_isRVC(alu_REG_0_isRVC)
  );
  UnpipelinedLSU lsu ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 57:19]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io__in_valid(lsu_io__in_valid),
    .io__in_bits_src1(lsu_io__in_bits_src1),
    .io__in_bits_src2(lsu_io__in_bits_src2),
    .io__in_bits_func(lsu_io__in_bits_func),
    .io__out_ready(lsu_io__out_ready),
    .io__out_valid(lsu_io__out_valid),
    .io__out_bits(lsu_io__out_bits),
    .io__wdata(lsu_io__wdata),
    .io__instr(lsu_io__instr),
    .io__dmem_req_ready(lsu_io__dmem_req_ready),
    .io__dmem_req_valid(lsu_io__dmem_req_valid),
    .io__dmem_req_bits_addr(lsu_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(lsu_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(lsu_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(lsu_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(lsu_io__dmem_req_bits_wdata),
    .io__dmem_resp_valid(lsu_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(lsu_io__dmem_resp_bits_rdata),
    .io__isMMIO(lsu_io__isMMIO),
    .io__dtlbPF(lsu_io__dtlbPF),
    .io__dtlbAF(lsu_io__dtlbAF),
    .io__vaddr(lsu_io__vaddr),
    .io__loadAddrMisaligned(lsu_io__loadAddrMisaligned),
    .io__storeAddrMisaligned(lsu_io__storeAddrMisaligned),
    .io__loadAccessFault(lsu_io__loadAccessFault),
    .io__storeAccessFault(lsu_io__storeAccessFault),
    .setLr_0(lsu_setLr_0),
    .lr_0(lsu_lr_0),
    .scInflight_0(lsu_scInflight_0),
    .amoReq_0(lsu_amoReq_0),
    .lr_addr(lsu_lr_addr),
    .dtlb_paddr(lsu_dtlb_paddr),
    ._T_12_0(lsu__T_12_0),
    .scIsSuccess_0(lsu_scIsSuccess_0),
    .setLrVal_0(lsu_setLrVal_0),
    .vmEnable(lsu_vmEnable),
    .DTLBFINISH(lsu_DTLBFINISH),
    .lsuMMIO_0(lsu_lsuMMIO_0),
    ._T_13_1(lsu__T_13_1),
    .setLrAddr_0(lsu_setLrAddr_0)
  );
  MDU mdu ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 66:19]
    .clock(mdu_clock),
    .reset(mdu_reset),
    .io_in_ready(mdu_io_in_ready),
    .io_in_valid(mdu_io_in_valid),
    .io_in_bits_src1(mdu_io_in_bits_src1),
    .io_in_bits_src2(mdu_io_in_bits_src2),
    .io_in_bits_func(mdu_io_in_bits_func),
    .io_out_ready(mdu_io_out_ready),
    .io_out_valid(mdu_io_out_valid),
    .io_out_bits(mdu_io_out_bits)
  );
  CSR csr ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 71:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_in_valid(csr_io_in_valid),
    .io_in_bits_src1(csr_io_in_bits_src1),
    .io_in_bits_src2(csr_io_in_bits_src2),
    .io_in_bits_func(csr_io_in_bits_func),
    .io_out_ready(csr_io_out_ready),
    .io_out_valid(csr_io_out_valid),
    .io_out_bits(csr_io_out_bits),
    .io_cfIn_instr(csr_io_cfIn_instr),
    .io_cfIn_pc(csr_io_cfIn_pc),
    .io_cfIn_exceptionVec_1(csr_io_cfIn_exceptionVec_1),
    .io_cfIn_exceptionVec_2(csr_io_cfIn_exceptionVec_2),
    .io_cfIn_exceptionVec_4(csr_io_cfIn_exceptionVec_4),
    .io_cfIn_exceptionVec_5(csr_io_cfIn_exceptionVec_5),
    .io_cfIn_exceptionVec_6(csr_io_cfIn_exceptionVec_6),
    .io_cfIn_exceptionVec_7(csr_io_cfIn_exceptionVec_7),
    .io_cfIn_exceptionVec_12(csr_io_cfIn_exceptionVec_12),
    .io_cfIn_exceptionVec_13(csr_io_cfIn_exceptionVec_13),
    .io_cfIn_exceptionVec_15(csr_io_cfIn_exceptionVec_15),
    .io_cfIn_intrVec_1(csr_io_cfIn_intrVec_1),
    .io_cfIn_intrVec_3(csr_io_cfIn_intrVec_3),
    .io_cfIn_intrVec_5(csr_io_cfIn_intrVec_5),
    .io_cfIn_intrVec_7(csr_io_cfIn_intrVec_7),
    .io_cfIn_intrVec_9(csr_io_cfIn_intrVec_9),
    .io_cfIn_intrVec_11(csr_io_cfIn_intrVec_11),
    .io_cfIn_crossBoundaryFault(csr_io_cfIn_crossBoundaryFault),
    .io_redirect_target(csr_io_redirect_target),
    .io_redirect_valid(csr_io_redirect_valid),
    .io_instrValid(csr_io_instrValid),
    .io_illegalJump_valid(csr_io_illegalJump_valid),
    .io_illegalJump_bits(csr_io_illegalJump_bits),
    .io_dmemExceptionAddr(csr_io_dmemExceptionAddr),
    .io_xretIsIllegal_ready(csr_io_xretIsIllegal_ready),
    .io_xretIsIllegal_valid(csr_io_xretIsIllegal_valid),
    .io_xretIsIllegal_bits(csr_io_xretIsIllegal_bits),
    .io_imemMMU_priviledgeMode(csr_io_imemMMU_priviledgeMode),
    .io_dmemMMU_priviledgeMode(csr_io_dmemMMU_priviledgeMode),
    .io_dmemMMU_status_sum(csr_io_dmemMMU_status_sum),
    .io_dmemMMU_status_mxr(csr_io_dmemMMU_status_mxr),
    .io_dmemMMU_loadPF(csr_io_dmemMMU_loadPF),
    .io_dmemMMU_storePF(csr_io_dmemMMU_storePF),
    .io_dmemMMU_laf(csr_io_dmemMMU_laf),
    .io_dmemMMU_saf(csr_io_dmemMMU_saf),
    .io_wenFix(csr_io_wenFix),
    .io_isPerfRead(csr_io_isPerfRead),
    .io_isExit(csr_io_isExit),
    .io_vmEnable(csr_io_vmEnable),
    .io_rfWenReal(csr_io_rfWenReal),
    .io_sfence_vma_invalid(csr_io_sfence_vma_invalid),
    .io_wfi_invalid(csr_io_wfi_invalid),
    .set_lr(csr_set_lr),
    .lr_0(csr_lr_0),
    .meip_0(csr_meip_0),
    .lrAddr_0(csr_lrAddr_0),
    .satp_0(csr_satp_0),
    .mtip_0(csr_mtip_0),
    .perfCntCondMultiCommit(csr_perfCntCondMultiCommit),
    .set_lr_val(csr_set_lr_val),
    .intrVecIDU_0(csr_intrVecIDU_0),
    .set_lr_addr(csr_set_lr_addr),
    .msip_0(csr_msip_0),
    .perfCntCondMinstret(csr_perfCntCondMinstret)
  );
  MOU mou ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 115:19]
    .clock(mou_clock),
    .reset(mou_reset),
    .io_in_valid(mou_io_in_valid),
    .io_in_bits_func(mou_io_in_bits_func),
    .io_cfIn_pc(mou_io_cfIn_pc),
    .io_redirect_target(mou_io_redirect_target),
    .io_redirect_valid(mou_io_redirect_valid),
    .flushICache_0(mou_flushICache_0),
    .flushTLB_0(mou_flushTLB_0)
  );
  EXUDiffWrapper diffMod ( // @[src/main/scala/nutcore/backend/seq/EXU.scala 170:25]
    .clock(diffMod_clock),
    .reset(diffMod_reset),
    .io_in_valid(diffMod_io_in_valid),
    .io_in_bits_cf_pc(diffMod_io_in_bits_cf_pc),
    .io_in_bits_ctrl_isNutCoreTrap(diffMod_io_in_bits_ctrl_isNutCoreTrap),
    .io_in_bits_data_src1(diffMod_io_in_bits_data_src1),
    .io_flush(diffMod_io_flush),
    .perfCntCondMinstret(diffMod_perfCntCondMinstret)
  );
  assign io__in_ready = ~io__in_valid | io__out_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 154:31]
  assign io__out_valid = io__in_valid & _io_out_valid_T_4; // @[src/main/scala/nutcore/backend/seq/EXU.scala 143:31]
  assign io__out_bits_decode_cf_instr = io__in_bits_cf_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 131:31]
  assign io__out_bits_decode_cf_pc = io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 130:28]
  assign io__out_bits_decode_cf_redirect_target = mou_io_redirect_valid ? mou_io_redirect_target :
    _io_out_bits_decode_cf_redirect_T_target; // @[src/main/scala/nutcore/backend/seq/EXU.scala 136:8]
  assign io__out_bits_decode_cf_redirect_valid = mou_io_redirect_valid ? mou_io_redirect_valid :
    _io_out_bits_decode_cf_redirect_T_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 136:8]
  assign io__out_bits_decode_ctrl_fuType = io__in_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/seq/EXU.scala 128:14]
  assign io__out_bits_decode_ctrl_rfWen = io__in_bits_ctrl_rfWen & (~hasException | ~fuValids_1) & ~(csr_io_wenFix &
    fuValids_3); // @[src/main/scala/nutcore/backend/seq/EXU.scala 126:68]
  assign io__out_bits_decode_ctrl_rfDest = io__in_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/seq/EXU.scala 127:14]
  assign io__out_bits_isMMIO = io__out_bits_decode_ctrl_rfWen & csr_io_isPerfRead | lsu_io__isMMIO; // @[src/main/scala/nutcore/backend/seq/EXU.scala 111:61 112:24 62:22]
  assign io__out_bits_commits_0 = alu_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 148:35]
  assign io__out_bits_commits_1 = lsu_io__out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 149:35]
  assign io__out_bits_commits_2 = mdu_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 151:35]
  assign io__out_bits_commits_3 = csr_io_out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 150:35]
  assign io__out_bits_isExit = csr_io_isExit; // @[src/main/scala/nutcore/backend/seq/EXU.scala 134:22]
  assign io__dmem_req_valid = lsu_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign io__dmem_req_bits_addr = lsu_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign io__dmem_req_bits_size = lsu_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign io__dmem_req_bits_cmd = lsu_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign io__dmem_req_bits_wmask = lsu_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign io__dmem_req_bits_wdata = lsu_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign io__forward_valid = io__in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 156:20]
  assign io__forward_wb_rfWen = io__in_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/seq/EXU.scala 157:23]
  assign io__forward_wb_rfDest = io__in_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/seq/EXU.scala 158:24]
  assign io__forward_wb_rfData = _io_forward_wb_rfData_T ? alu_io_out_bits : lsu_io__out_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 159:30]
  assign io__forward_fuType = io__in_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/seq/EXU.scala 160:21]
  assign io__memMMU_imem_priviledgeMode = csr_io_imemMMU_priviledgeMode; // @[src/main/scala/nutcore/backend/seq/EXU.scala 89:18]
  assign io__memMMU_dmem_priviledgeMode = csr_io_dmemMMU_priviledgeMode; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign io__memMMU_dmem_status_sum = csr_io_dmemMMU_status_sum; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign io__memMMU_dmem_status_mxr = csr_io_dmemMMU_status_mxr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign io__sfence_vma_invalid = csr_io_sfence_vma_invalid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 86:25]
  assign io__wfi_invalid = csr_io_wfi_invalid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 87:18]
  assign lr = csr_lr_0;
  assign scInflight = lsu_scInflight_0;
  assign REG_valid = alu_REG_0_valid;
  assign REG_pc = alu_REG_0_pc;
  assign REG_isMissPredict = alu_REG_0_isMissPredict;
  assign REG_actualTarget = alu_REG_0_actualTarget;
  assign REG_fuOpType = alu_REG_0_fuOpType;
  assign REG_btbType = alu_REG_0_btbType;
  assign REG_isRVC = alu_REG_0_isRVC;
  assign amoReq = lsu_amoReq_0;
  assign lrAddr = csr_lrAddr_0;
  assign satp = csr_satp_0;
  assign flushICache = mou_flushICache_0;
  assign flushTLB = mou_flushTLB_0;
  assign intrVecIDU = csr_intrVecIDU_0;
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_in_valid = _T | _T_1 ? 1'h0 : io__in_bits_ctrl_fuType == 3'h0 & io__in_valid & ~io__flush & ~(|
    _fuValids_0_T_4); // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  assign alu_io_in_bits_src1 = io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 41:34]
  assign alu_io_in_bits_src2 = io__in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 42:34]
  assign alu_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/ALU.scala 85:15]
  assign alu_io_out_ready = 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 53:20]
  assign alu_io_cfIn_instr = io__in_bits_cf_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 51:15]
  assign alu_io_cfIn_pc = io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 51:15]
  assign alu_io_cfIn_pnpc = io__in_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 51:15]
  assign alu_io_cfIn_brIdx = io__in_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/seq/EXU.scala 51:15]
  assign alu_io_offset = io__in_bits_data_imm; // @[src/main/scala/nutcore/backend/seq/EXU.scala 52:17]
  assign alu_io_iVmEnable = csr_io_vmEnable; // @[src/main/scala/nutcore/backend/seq/EXU.scala 90:20]
  assign alu_io_jumpIsIllegal_ready = io__in_valid & _fuValids_0_T_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 97:45]
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io__in_valid = _T | _T_1 ? 1'h0 : io__in_bits_ctrl_fuType == 3'h1 & io__in_valid & ~io__flush & ~(|
    _fuValids_0_T_4); // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  assign lsu_io__in_bits_src1 = io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 41:34]
  assign lsu_io__in_bits_src2 = io__in_bits_data_imm; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 51:21]
  assign lsu_io__in_bits_func = io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/UnpipelinedLSU.scala 52:21]
  assign lsu_io__out_ready = 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 64:20]
  assign lsu_io__wdata = io__in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 42:34]
  assign lsu_io__instr = io__in_bits_cf_instr[31:0]; // @[src/main/scala/nutcore/backend/seq/EXU.scala 61:16]
  assign lsu_io__dmem_req_ready = io__dmem_req_ready; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign lsu_io__dmem_resp_valid = io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign lsu_io__dmem_resp_bits_rdata = io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/seq/EXU.scala 63:11]
  assign lsu_lr_0 = lr;
  assign lsu_lr_addr = lrAddr;
  assign lsu_dtlb_paddr = paddr;
  assign lsu__T_12_0 = _T_12_0;
  assign lsu_scIsSuccess_0 = scIsSuccess;
  assign lsu_vmEnable = vmEnable;
  assign lsu_DTLBFINISH = tlbFinish;
  assign lsu_lsuMMIO_0 = ismmio;
  assign lsu__T_13_1 = _T_13_1;
  assign mdu_clock = clock;
  assign mdu_reset = reset;
  assign mdu_io_in_valid = _T | _T_1 ? 1'h0 : io__in_bits_ctrl_fuType == 3'h2 & io__in_valid & ~io__flush & ~(|
    _fuValids_0_T_4); // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  assign mdu_io_in_bits_src1 = io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 41:34]
  assign mdu_io_in_bits_src2 = io__in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 42:34]
  assign mdu_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/MDU.scala 143:15]
  assign mdu_io_out_ready = 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 68:20]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_in_valid = _T | _T_1 | io__in_bits_ctrl_fuType == 3'h3 & io__in_valid & ~io__flush & ~(|_fuValids_0_T_4)
    ; // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  assign csr_io_in_bits_src1 = io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 41:34]
  assign csr_io_in_bits_src2 = io__in_bits_data_src2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 42:34]
  assign csr_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/CSR.scala 207:15]
  assign csr_io_out_ready = 1'h1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 84:20]
  assign csr_io_cfIn_instr = io__in_bits_cf_instr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_pc = io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_exceptionVec_1 = _T | _T_1 ? _GEN_1 : io__in_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15 99:65]
  assign csr_io_cfIn_exceptionVec_2 = io__in_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_exceptionVec_4 = lsu_io__loadAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 74:48]
  assign csr_io_cfIn_exceptionVec_5 = lsu_io__loadAccessFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 76:45]
  assign csr_io_cfIn_exceptionVec_6 = lsu_io__storeAddrMisaligned; // @[src/main/scala/nutcore/backend/seq/EXU.scala 75:49]
  assign csr_io_cfIn_exceptionVec_7 = lsu_io__storeAccessFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 77:46]
  assign csr_io_cfIn_exceptionVec_12 = _T | _T_1 ? _GEN_0 : io__in_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15 99:65]
  assign csr_io_cfIn_exceptionVec_13 = lsu_io__in_valid & lsu_io__dtlbPF & _csr_io_cfIn_exceptionVec_13_T_7; // @[src/main/scala/nutcore/backend/seq/EXU.scala 78:79]
  assign csr_io_cfIn_exceptionVec_15 = _csr_io_cfIn_exceptionVec_13_T & _csr_io_cfIn_exceptionVec_13_T_6; // @[src/main/scala/nutcore/backend/seq/EXU.scala 79:80]
  assign csr_io_cfIn_intrVec_1 = io__in_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_intrVec_3 = io__in_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_intrVec_5 = io__in_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_intrVec_7 = io__in_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_intrVec_9 = io__in_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_intrVec_11 = io__in_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_cfIn_crossBoundaryFault = io__in_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/backend/seq/EXU.scala 73:15]
  assign csr_io_instrValid = io__in_valid & _fuValids_0_T_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 80:36]
  assign csr_io_illegalJump_valid = alu_io_jumpIsIllegal_valid | csr_io_xretIsIllegal_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 95:60]
  assign csr_io_illegalJump_bits = alu_io_jumpIsIllegal_valid ? alu_io_jumpIsIllegal_bits : csr_io_xretIsIllegal_bits; // @[src/main/scala/nutcore/backend/seq/EXU.scala 96:36]
  assign csr_io_dmemExceptionAddr = lsu_io__vaddr; // @[src/main/scala/nutcore/backend/seq/EXU.scala 92:28]
  assign csr_io_xretIsIllegal_ready = io__in_valid & _fuValids_0_T_2; // @[src/main/scala/nutcore/backend/seq/EXU.scala 98:45]
  assign csr_io_dmemMMU_loadPF = io__memMMU_dmem_loadPF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign csr_io_dmemMMU_storePF = io__memMMU_dmem_storePF; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign csr_io_dmemMMU_laf = io__memMMU_dmem_laf; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign csr_io_dmemMMU_saf = io__memMMU_dmem_saf; // @[src/main/scala/nutcore/backend/seq/EXU.scala 91:18]
  assign csr_io_rfWenReal = io__in_bits_ctrl_rfWen & io__in_bits_ctrl_rfDest != 5'h0; // @[src/main/scala/nutcore/backend/seq/EXU.scala 85:45]
  assign csr_set_lr = lsu_setLr_0;
  assign csr_meip_0 = io_extra_meip_0;
  assign csr_mtip_0 = io_extra_mtip;
  assign csr_perfCntCondMultiCommit = falseWire;
  assign csr_set_lr_val = lsu_setLrVal_0;
  assign csr_set_lr_addr = lsu_setLrAddr_0;
  assign csr_msip_0 = io_extra_msip;
  assign csr_perfCntCondMinstret = io_in_valid;
  assign mou_clock = clock;
  assign mou_reset = reset;
  assign mou_io_in_valid = _T | _T_1 ? 1'h0 : io__in_bits_ctrl_fuType == 3'h4 & io__in_valid & ~io__flush & ~(|
    _fuValids_0_T_4); // @[src/main/scala/nutcore/backend/seq/EXU.scala 99:65 101:9 47:46]
  assign mou_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/fu/MOU.scala 45:15]
  assign mou_io_cfIn_pc = io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 118:15]
  assign diffMod_clock = clock;
  assign diffMod_reset = reset;
  assign diffMod_io_in_valid = io__in_valid; // @[src/main/scala/nutcore/backend/seq/EXU.scala 171:25]
  assign diffMod_io_in_bits_cf_pc = io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/seq/EXU.scala 172:24]
  assign diffMod_io_in_bits_ctrl_isNutCoreTrap = io__in_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/seq/EXU.scala 172:24]
  assign diffMod_io_in_bits_data_src1 = io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/seq/EXU.scala 172:24]
  assign diffMod_io_flush = io__flush; // @[src/main/scala/nutcore/backend/seq/EXU.scala 173:22]
  assign diffMod_perfCntCondMinstret = io_in_valid;
endmodule
module DummyDPICWrapper_4(
  input         clock,
  input         reset,
  input         io_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_skip, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_isRVC, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_rfwen, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [4:0]  io_bits_wpdest, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [7:0]  io_bits_wdest, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_pc, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [31:0] io_bits_instr, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [7:0]  io_bits_special // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_valid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_skip; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_isRVC; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_rfwen; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_fpwen; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_vecwen; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [4:0] dpic_io_wpdest; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_wdest; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_pc; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [31:0] dpic_io_instr; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [9:0] dpic_io_robIdx; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [6:0] dpic_io_lqIdx; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [6:0] dpic_io_sqIdx; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_isLoad; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_isStore; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_nFused; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_special; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_index; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestInstrCommit dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_valid(dpic_io_valid),
    .io_skip(dpic_io_skip),
    .io_isRVC(dpic_io_isRVC),
    .io_rfwen(dpic_io_rfwen),
    .io_fpwen(dpic_io_fpwen),
    .io_vecwen(dpic_io_vecwen),
    .io_wpdest(dpic_io_wpdest),
    .io_wdest(dpic_io_wdest),
    .io_pc(dpic_io_pc),
    .io_instr(dpic_io_instr),
    .io_robIdx(dpic_io_robIdx),
    .io_lqIdx(dpic_io_lqIdx),
    .io_sqIdx(dpic_io_sqIdx),
    .io_isLoad(dpic_io_isLoad),
    .io_isStore(dpic_io_isStore),
    .io_nFused(dpic_io_nFused),
    .io_special(dpic_io_special),
    .io_coreid(dpic_io_coreid),
    .io_index(dpic_io_index)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = io_valid; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_valid = io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_skip = io_bits_skip; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_isRVC = io_bits_isRVC; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_rfwen = io_bits_rfwen; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_fpwen = 1'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_vecwen = 1'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_wpdest = io_bits_wpdest; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_wdest = io_bits_wdest; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_pc = io_bits_pc; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_instr = io_bits_instr; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_robIdx = 10'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_lqIdx = 7'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_sqIdx = 7'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_isLoad = 1'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_isStore = 1'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_nFused = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_special = io_bits_special; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_index = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module DiffInstrCommitWrapper(
  input         clock,
  input         reset,
  input         io_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 68:18]
  input         io_skip, // @[src/main/scala/nutcore/backend/seq/WBU.scala 68:18]
  input         io_isRVC, // @[src/main/scala/nutcore/backend/seq/WBU.scala 68:18]
  input         io_rfwen, // @[src/main/scala/nutcore/backend/seq/WBU.scala 68:18]
  input  [4:0]  io_wpdest, // @[src/main/scala/nutcore/backend/seq/WBU.scala 68:18]
  input  [7:0]  io_wdest, // @[src/main/scala/nutcore/backend/seq/WBU.scala 68:18]
  input  [63:0] io_pc, // @[src/main/scala/nutcore/backend/seq/WBU.scala 68:18]
  input  [31:0] io_instr, // @[src/main/scala/nutcore/backend/seq/WBU.scala 68:18]
  input  [7:0]  io_special // @[src/main/scala/nutcore/backend/seq/WBU.scala 68:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  difftest_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_skip; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_isRVC; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_rfwen; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [4:0] difftest_module_io_bits_wpdest; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [7:0] difftest_module_io_bits_wdest; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_pc; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [31:0] difftest_module_io_bits_instr; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [7:0] difftest_module_io_bits_special; // @[difftest/src/main/scala/DPIC.scala 299:24]
  reg  difftest_REG_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
  reg  difftest_REG_skip; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
  reg  difftest_REG_isRVC; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
  reg  difftest_REG_rfwen; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
  reg [4:0] difftest_REG_wpdest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
  reg [7:0] difftest_REG_wdest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
  reg [63:0] difftest_REG_pc; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
  reg [31:0] difftest_REG_instr; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
  reg [7:0] difftest_REG_special; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
  DummyDPICWrapper_4 difftest_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_clock),
    .reset(difftest_module_reset),
    .io_valid(difftest_module_io_valid),
    .io_bits_valid(difftest_module_io_bits_valid),
    .io_bits_skip(difftest_module_io_bits_skip),
    .io_bits_isRVC(difftest_module_io_bits_isRVC),
    .io_bits_rfwen(difftest_module_io_bits_rfwen),
    .io_bits_wpdest(difftest_module_io_bits_wpdest),
    .io_bits_wdest(difftest_module_io_bits_wdest),
    .io_bits_pc(difftest_module_io_bits_pc),
    .io_bits_instr(difftest_module_io_bits_instr),
    .io_bits_special(difftest_module_io_bits_special)
  );
  assign difftest_module_clock = clock;
  assign difftest_module_reset = reset;
  assign difftest_module_io_valid = difftest_REG_valid; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 71:16]
  assign difftest_module_io_bits_valid = difftest_REG_valid; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 71:16]
  assign difftest_module_io_bits_skip = difftest_REG_skip; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 71:16]
  assign difftest_module_io_bits_isRVC = difftest_REG_isRVC; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 71:16]
  assign difftest_module_io_bits_rfwen = difftest_REG_rfwen; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 71:16]
  assign difftest_module_io_bits_wpdest = difftest_REG_wpdest; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 71:16]
  assign difftest_module_io_bits_wdest = difftest_REG_wdest; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 71:16]
  assign difftest_module_io_bits_pc = difftest_REG_pc; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 71:16]
  assign difftest_module_io_bits_instr = difftest_REG_instr; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 71:16]
  assign difftest_module_io_bits_special = difftest_REG_special; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 71:16]
  always @(posedge clock) begin
    difftest_REG_valid <= io_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
    difftest_REG_skip <= io_skip; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
    difftest_REG_isRVC <= io_isRVC; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
    difftest_REG_rfwen <= io_rfwen; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
    difftest_REG_wpdest <= io_wpdest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
    difftest_REG_wdest <= io_wdest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
    difftest_REG_pc <= io_pc; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
    difftest_REG_instr <= io_instr; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
    difftest_REG_special <= io_special; // @[src/main/scala/nutcore/backend/seq/WBU.scala 71:26]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  difftest_REG_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  difftest_REG_skip = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  difftest_REG_isRVC = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  difftest_REG_rfwen = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  difftest_REG_wpdest = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  difftest_REG_wdest = _RAND_5[7:0];
  _RAND_6 = {2{`RANDOM}};
  difftest_REG_pc = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  difftest_REG_instr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  difftest_REG_special = _RAND_8[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DummyDPICWrapper_5(
  input         clock,
  input         reset,
  input         io_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input         io_bits_valid, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [4:0]  io_bits_address, // @[difftest/src/main/scala/DPIC.scala 272:14]
  input  [63:0] io_bits_data // @[difftest/src/main/scala/DPIC.scala 272:14]
);
  wire  dpic_clock; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_enable; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire  dpic_io_valid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [4:0] dpic_io_address; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [63:0] dpic_io_data; // @[difftest/src/main/scala/DPIC.scala 273:20]
  wire [7:0] dpic_io_coreid; // @[difftest/src/main/scala/DPIC.scala 273:20]
  DifftestIntWriteback dpic ( // @[difftest/src/main/scala/DPIC.scala 273:20]
    .clock(dpic_clock),
    .enable(dpic_enable),
    .io_valid(dpic_io_valid),
    .io_address(dpic_io_address),
    .io_data(dpic_io_data),
    .io_coreid(dpic_io_coreid)
  );
  assign dpic_clock = clock; // @[difftest/src/main/scala/DPIC.scala 274:14]
  assign dpic_enable = io_valid; // @[difftest/src/main/scala/DPIC.scala 275:27]
  assign dpic_io_valid = io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_address = io_bits_address; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_data = io_bits_data; // @[difftest/src/main/scala/DPIC.scala 277:11]
  assign dpic_io_coreid = 8'h0; // @[difftest/src/main/scala/DPIC.scala 277:11]
endmodule
module DiffIntWbWrapper(
  input         clock,
  input         reset,
  input         io_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 104:18]
  input  [4:0]  io_address, // @[src/main/scala/nutcore/backend/seq/WBU.scala 104:18]
  input  [63:0] io_data // @[src/main/scala/nutcore/backend/seq/WBU.scala 104:18]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  difftest_module_clock; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_reset; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire  difftest_module_io_bits_valid; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [4:0] difftest_module_io_bits_address; // @[difftest/src/main/scala/DPIC.scala 299:24]
  wire [63:0] difftest_module_io_bits_data; // @[difftest/src/main/scala/DPIC.scala 299:24]
  reg  difftest_REG_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 106:26]
  reg [4:0] difftest_REG_address; // @[src/main/scala/nutcore/backend/seq/WBU.scala 106:26]
  reg [63:0] difftest_REG_data; // @[src/main/scala/nutcore/backend/seq/WBU.scala 106:26]
  DummyDPICWrapper_5 difftest_module ( // @[difftest/src/main/scala/DPIC.scala 299:24]
    .clock(difftest_module_clock),
    .reset(difftest_module_reset),
    .io_valid(difftest_module_io_valid),
    .io_bits_valid(difftest_module_io_bits_valid),
    .io_bits_address(difftest_module_io_bits_address),
    .io_bits_data(difftest_module_io_bits_data)
  );
  assign difftest_module_clock = clock;
  assign difftest_module_reset = reset;
  assign difftest_module_io_valid = difftest_REG_valid; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 106:16]
  assign difftest_module_io_bits_valid = difftest_REG_valid; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 106:16]
  assign difftest_module_io_bits_address = difftest_REG_address; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 106:16]
  assign difftest_module_io_bits_data = difftest_REG_data; // @[difftest/src/main/scala/Difftest.scala 460:27 src/main/scala/nutcore/backend/seq/WBU.scala 106:16]
  always @(posedge clock) begin
    difftest_REG_valid <= io_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 106:26]
    difftest_REG_address <= io_address; // @[src/main/scala/nutcore/backend/seq/WBU.scala 106:26]
    difftest_REG_data <= io_data; // @[src/main/scala/nutcore/backend/seq/WBU.scala 106:26]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  difftest_REG_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  difftest_REG_address = _RAND_1[4:0];
  _RAND_2 = {2{`RANDOM}};
  difftest_REG_data = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WBU(
  input         clock,
  input         reset,
  input         io__in_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_decode_cf_instr, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [38:0] io__in_bits_decode_cf_pc, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [38:0] io__in_bits_decode_cf_redirect_target, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input         io__in_bits_decode_cf_redirect_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [2:0]  io__in_bits_decode_ctrl_fuType, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input         io__in_bits_decode_ctrl_rfWen, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [4:0]  io__in_bits_decode_ctrl_rfDest, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input         io__in_bits_isMMIO, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_commits_0, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_commits_1, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_commits_2, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input  [63:0] io__in_bits_commits_3, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  input         io__in_bits_isExit, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output        io__wb_rfWen, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output [4:0]  io__wb_rfDest, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output [63:0] io__wb_rfData, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output [38:0] io__redirect_target, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output        io__redirect_valid, // @[src/main/scala/nutcore/backend/seq/WBU.scala 29:14]
  output        falseWire_0,
  output        io_in_valid
);
  wire  DiffInstrCommitWrapper_clock; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire  DiffInstrCommitWrapper_reset; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire  DiffInstrCommitWrapper_io_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire  DiffInstrCommitWrapper_io_skip; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire  DiffInstrCommitWrapper_io_isRVC; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire  DiffInstrCommitWrapper_io_rfwen; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire [4:0] DiffInstrCommitWrapper_io_wpdest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire [7:0] DiffInstrCommitWrapper_io_wdest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire [63:0] DiffInstrCommitWrapper_io_pc; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire [31:0] DiffInstrCommitWrapper_io_instr; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire [7:0] DiffInstrCommitWrapper_io_special; // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
  wire  DiffIntWbWrapper_clock; // @[src/main/scala/nutcore/backend/seq/WBU.scala 114:26]
  wire  DiffIntWbWrapper_reset; // @[src/main/scala/nutcore/backend/seq/WBU.scala 114:26]
  wire  DiffIntWbWrapper_io_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 114:26]
  wire [4:0] DiffIntWbWrapper_io_address; // @[src/main/scala/nutcore/backend/seq/WBU.scala 114:26]
  wire [63:0] DiffIntWbWrapper_io_data; // @[src/main/scala/nutcore/backend/seq/WBU.scala 114:26]
  wire [63:0] _GEN_1 = 3'h1 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_1 : io__in_bits_commits_0; // @[src/main/scala/nutcore/backend/seq/WBU.scala 37:{16,16}]
  wire [63:0] _GEN_2 = 3'h2 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_2 : _GEN_1; // @[src/main/scala/nutcore/backend/seq/WBU.scala 37:{16,16}]
  wire [63:0] _GEN_3 = 3'h3 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_3 : _GEN_2; // @[src/main/scala/nutcore/backend/seq/WBU.scala 37:{16,16}]
  wire  signBit = io__in_bits_decode_cf_pc[38]; // @[src/main/scala/utils/BitUtils.scala 41:20]
  wire [24:0] _T = signBit ? 25'h1ffffff : 25'h0; // @[src/main/scala/utils/BitUtils.scala 42:46]
  wire  _T_4 = io__wb_rfDest != 5'h0; // @[src/main/scala/nutcore/backend/seq/WBU.scala 89:51]
  wire [1:0] _T_6 = {io__in_bits_isExit,1'h0}; // @[difftest/src/main/scala/Bundles.scala 81:19]
  wire  falseWire = 1'h0; // @[src/main/scala/nutcore/backend/seq/WBU.scala 62:{27,27}]
  DiffInstrCommitWrapper DiffInstrCommitWrapper ( // @[src/main/scala/nutcore/backend/seq/WBU.scala 82:26]
    .clock(DiffInstrCommitWrapper_clock),
    .reset(DiffInstrCommitWrapper_reset),
    .io_valid(DiffInstrCommitWrapper_io_valid),
    .io_skip(DiffInstrCommitWrapper_io_skip),
    .io_isRVC(DiffInstrCommitWrapper_io_isRVC),
    .io_rfwen(DiffInstrCommitWrapper_io_rfwen),
    .io_wpdest(DiffInstrCommitWrapper_io_wpdest),
    .io_wdest(DiffInstrCommitWrapper_io_wdest),
    .io_pc(DiffInstrCommitWrapper_io_pc),
    .io_instr(DiffInstrCommitWrapper_io_instr),
    .io_special(DiffInstrCommitWrapper_io_special)
  );
  DiffIntWbWrapper DiffIntWbWrapper ( // @[src/main/scala/nutcore/backend/seq/WBU.scala 114:26]
    .clock(DiffIntWbWrapper_clock),
    .reset(DiffIntWbWrapper_reset),
    .io_valid(DiffIntWbWrapper_io_valid),
    .io_address(DiffIntWbWrapper_io_address),
    .io_data(DiffIntWbWrapper_io_data)
  );
  assign io__wb_rfWen = io__in_bits_decode_ctrl_rfWen & io__in_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 35:47]
  assign io__wb_rfDest = io__in_bits_decode_ctrl_rfDest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 36:16]
  assign io__wb_rfData = 3'h4 == io__in_bits_decode_ctrl_fuType ? 64'h0 : _GEN_3; // @[src/main/scala/nutcore/backend/seq/WBU.scala 37:{16,16}]
  assign io__redirect_target = io__in_bits_decode_cf_redirect_target; // @[src/main/scala/nutcore/backend/seq/WBU.scala 41:15]
  assign io__redirect_valid = io__in_bits_decode_cf_redirect_valid & io__in_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 42:60]
  assign falseWire_0 = falseWire;
  assign io_in_valid = io__in_valid;
  assign DiffInstrCommitWrapper_clock = clock;
  assign DiffInstrCommitWrapper_reset = reset;
  assign DiffInstrCommitWrapper_io_valid = io__in_valid; // @[src/main/scala/nutcore/backend/seq/WBU.scala 84:20]
  assign DiffInstrCommitWrapper_io_skip = io__in_bits_isMMIO; // @[src/main/scala/nutcore/backend/seq/WBU.scala 87:19]
  assign DiffInstrCommitWrapper_io_isRVC = io__in_bits_decode_cf_instr[1:0] != 2'h3; // @[src/main/scala/nutcore/backend/seq/WBU.scala 88:56]
  assign DiffInstrCommitWrapper_io_rfwen = io__wb_rfWen & io__wb_rfDest != 5'h0; // @[src/main/scala/nutcore/backend/seq/WBU.scala 89:35]
  assign DiffInstrCommitWrapper_io_wpdest = io__wb_rfDest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 91:21]
  assign DiffInstrCommitWrapper_io_wdest = {{3'd0}, io__wb_rfDest}; // @[src/main/scala/nutcore/backend/seq/WBU.scala 90:20]
  assign DiffInstrCommitWrapper_io_pc = {_T,io__in_bits_decode_cf_pc}; // @[src/main/scala/utils/BitUtils.scala 42:41]
  assign DiffInstrCommitWrapper_io_instr = io__in_bits_decode_cf_instr[31:0]; // @[src/main/scala/nutcore/backend/seq/WBU.scala 86:20]
  assign DiffInstrCommitWrapper_io_special = {{6'd0}, _T_6}; // @[difftest/src/main/scala/Bundles.scala 81:13]
  assign DiffIntWbWrapper_clock = clock;
  assign DiffIntWbWrapper_reset = reset;
  assign DiffIntWbWrapper_io_valid = io__wb_rfWen & _T_4; // @[src/main/scala/nutcore/backend/seq/WBU.scala 116:35]
  assign DiffIntWbWrapper_io_address = io__wb_rfDest; // @[src/main/scala/nutcore/backend/seq/WBU.scala 117:22]
  assign DiffIntWbWrapper_io_data = io__wb_rfData; // @[src/main/scala/nutcore/backend/seq/WBU.scala 118:19]
endmodule
module Backend_inorder(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_valid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [63:0] io_in_0_bits_cf_instr, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [38:0] io_in_0_bits_cf_pc, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [38:0] io_in_0_bits_cf_pnpc, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_exceptionVec_1, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_exceptionVec_2, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_exceptionVec_12, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_1, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_3, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_5, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_7, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_9, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_intrVec_11, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [3:0]  io_in_0_bits_cf_brIdx, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_cf_crossBoundaryFault, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_ctrl_src1Type, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_ctrl_src2Type, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [2:0]  io_in_0_bits_ctrl_fuType, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [6:0]  io_in_0_bits_ctrl_fuOpType, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [4:0]  io_in_0_bits_ctrl_rfSrc1, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [4:0]  io_in_0_bits_ctrl_rfSrc2, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_ctrl_rfWen, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [4:0]  io_in_0_bits_ctrl_rfDest, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_in_0_bits_ctrl_isNutCoreTrap, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [63:0] io_in_0_bits_data_imm, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [1:0]  io_flush, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_dmem_req_ready, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_dmem_req_valid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [38:0] io_dmem_req_bits_addr, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [2:0]  io_dmem_req_bits_size, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [3:0]  io_dmem_req_bits_cmd, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [7:0]  io_dmem_req_bits_wmask, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [63:0] io_dmem_req_bits_wdata, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_dmem_resp_valid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input  [63:0] io_dmem_resp_bits_rdata, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [1:0]  io_memMMU_imem_priviledgeMode, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [1:0]  io_memMMU_dmem_priviledgeMode, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_memMMU_dmem_status_sum, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_memMMU_dmem_status_mxr, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_memMMU_dmem_loadPF, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_memMMU_dmem_storePF, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_memMMU_dmem_laf, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  input         io_memMMU_dmem_saf, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_sfence_vma_invalid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_wfi_invalid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output [38:0] io_redirect_target, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        io_redirect_valid, // @[src/main/scala/nutcore/backend/ooo/Backend.scala 669:14]
  output        lr,
  input         io_extra_meip_0,
  output        scInflight,
  output        REG_valid,
  output [38:0] REG_pc,
  output        REG_isMissPredict,
  output [38:0] REG_actualTarget,
  output [6:0]  REG_fuOpType,
  output [1:0]  REG_btbType,
  output        REG_isRVC,
  output        amoReq,
  output [63:0] lrAddr,
  input  [55:0] paddr,
  output [63:0] satp,
  input         _T_12,
  input         scIsSuccess,
  input         io_extra_mtip,
  output        flushICache,
  input         vmEnable,
  output        flushTLB,
  output [11:0] intrVecIDU,
  input         tlbFinish,
  input         ismmio,
  input         _T_13_0,
  input         io_extra_msip
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
`endif // RANDOMIZE_REG_INIT
  wire  isu_clock; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_reset; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_in_0_bits_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [38:0] isu_io_in_0_bits_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [38:0] isu_io_in_0_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [3:0] isu_io_in_0_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [2:0] isu_io_in_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [6:0] isu_io_in_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_in_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_in_0_bits_data_imm; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_out_bits_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [38:0] isu_io_out_bits_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [38:0] isu_io_out_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [3:0] isu_io_out_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [2:0] isu_io_out_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [6:0] isu_io_out_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] isu_io_out_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_out_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_out_bits_data_src1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_out_bits_data_src2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_out_bits_data_imm; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] isu_io_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_forward_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_forward_wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [4:0] isu_io_forward_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [63:0] isu_io_forward_wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire [2:0] isu_io_forward_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  isu_io_flush; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
  wire  exu_clock; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_reset; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__in_bits_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_io__in_bits_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_io__in_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [3:0] exu_io__in_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [2:0] exu_io__in_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [6:0] exu_io__in_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [4:0] exu_io__in_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__in_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__in_bits_data_src1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__in_bits_data_src2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__in_bits_data_imm; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__out_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__out_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__out_bits_decode_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_io__out_bits_decode_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_io__out_bits_decode_cf_redirect_target; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__out_bits_decode_cf_redirect_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [2:0] exu_io__out_bits_decode_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__out_bits_decode_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [4:0] exu_io__out_bits_decode_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__out_bits_isMMIO; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__out_bits_commits_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__out_bits_commits_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__out_bits_commits_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__out_bits_commits_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__out_bits_isExit; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__flush; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__dmem_req_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [2:0] exu_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [3:0] exu_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [7:0] exu_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__dmem_resp_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__forward_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__forward_wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [4:0] exu_io__forward_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_io__forward_wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [2:0] exu_io__forward_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [1:0] exu_io__memMMU_imem_priviledgeMode; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [1:0] exu_io__memMMU_dmem_priviledgeMode; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__memMMU_dmem_status_sum; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__memMMU_dmem_status_mxr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__memMMU_dmem_loadPF; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__memMMU_dmem_storePF; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__memMMU_dmem_laf; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__memMMU_dmem_saf; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__sfence_vma_invalid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io__wfi_invalid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_lr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io_extra_meip_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_scInflight; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_REG_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_REG_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_REG_isMissPredict; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [38:0] exu_REG_actualTarget; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [6:0] exu_REG_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [1:0] exu_REG_btbType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_REG_isRVC; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_amoReq; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_lrAddr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [55:0] exu_paddr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [63:0] exu_satp; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu__T_12_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_scIsSuccess; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io_extra_mtip; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_flushICache; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_falseWire; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_vmEnable; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_flushTLB; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire [11:0] exu_intrVecIDU; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_tlbFinish; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_ismmio; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu__T_13_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io_extra_msip; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  exu_io_in_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
  wire  wbu_clock; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_reset; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__in_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] wbu_io__in_bits_decode_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [38:0] wbu_io__in_bits_decode_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [38:0] wbu_io__in_bits_decode_cf_redirect_target; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__in_bits_decode_cf_redirect_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [2:0] wbu_io__in_bits_decode_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__in_bits_decode_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [4:0] wbu_io__in_bits_decode_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__in_bits_isMMIO; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] wbu_io__in_bits_commits_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] wbu_io__in_bits_commits_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] wbu_io__in_bits_commits_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] wbu_io__in_bits_commits_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__in_bits_isExit; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [4:0] wbu_io__wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [63:0] wbu_io__wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire [38:0] wbu_io__redirect_target; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io__redirect_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_falseWire_0; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  wbu_io_in_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
  wire  _T = exu_io__out_ready & exu_io__out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  valid; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _GEN_0 = _T ? 1'h0 : valid; // @[src/main/scala/utils/Pipeline.scala 24:24 25:{25,33}]
  wire  _T_2 = isu_io_out_valid & exu_io__in_ready; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  _GEN_1 = isu_io_out_valid & exu_io__in_ready | _GEN_0; // @[src/main/scala/utils/Pipeline.scala 26:{38,46}]
  reg [63:0] exu_io_in_bits_r_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] exu_io_in_bits_r_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] exu_io_in_bits_r_cf_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_exceptionVec_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_5; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_7; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_9; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_intrVec_11; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] exu_io_in_bits_r_cf_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_cf_crossBoundaryFault; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [2:0] exu_io_in_bits_r_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [6:0] exu_io_in_bits_r_ctrl_fuOpType; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [4:0] exu_io_in_bits_r_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  exu_io_in_bits_r_ctrl_isNutCoreTrap; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] exu_io_in_bits_r_data_src1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] exu_io_in_bits_r_data_src2; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] exu_io_in_bits_r_data_imm; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _T_4 = exu_io__out_valid; // @[src/main/scala/utils/Pipeline.scala 26:22]
  reg [63:0] wbu_io_in_bits_r_decode_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] wbu_io_in_bits_r_decode_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [38:0] wbu_io_in_bits_r_decode_cf_redirect_target; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  wbu_io_in_bits_r_decode_cf_redirect_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [2:0] wbu_io_in_bits_r_decode_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  wbu_io_in_bits_r_decode_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [4:0] wbu_io_in_bits_r_decode_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  wbu_io_in_bits_r_isMMIO; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_commits_0; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_commits_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_commits_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] wbu_io_in_bits_r_commits_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  wbu_io_in_bits_r_isExit; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  valid_p; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  valid_t = valid ^ valid_p; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  toggle_5404_clock;
  wire  toggle_5404_reset;
  wire  toggle_5404_valid;
  reg  toggle_5404_valid_reg;
  reg [63:0] exu_io_in_bits_r_cf_instr_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [63:0] exu_io_in_bits_r_cf_instr_t = exu_io_in_bits_r_cf_instr ^ exu_io_in_bits_r_cf_instr_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5405_clock;
  wire  toggle_5405_reset;
  wire [63:0] toggle_5405_valid;
  reg [63:0] toggle_5405_valid_reg;
  reg [38:0] exu_io_in_bits_r_cf_pc_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [38:0] exu_io_in_bits_r_cf_pc_t = exu_io_in_bits_r_cf_pc ^ exu_io_in_bits_r_cf_pc_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5469_clock;
  wire  toggle_5469_reset;
  wire [38:0] toggle_5469_valid;
  reg [38:0] toggle_5469_valid_reg;
  reg [38:0] exu_io_in_bits_r_cf_pnpc_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [38:0] exu_io_in_bits_r_cf_pnpc_t = exu_io_in_bits_r_cf_pnpc ^ exu_io_in_bits_r_cf_pnpc_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5508_clock;
  wire  toggle_5508_reset;
  wire [38:0] toggle_5508_valid;
  reg [38:0] toggle_5508_valid_reg;
  reg  exu_io_in_bits_r_cf_exceptionVec_1_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  exu_io_in_bits_r_cf_exceptionVec_1_t = exu_io_in_bits_r_cf_exceptionVec_1 ^ exu_io_in_bits_r_cf_exceptionVec_1_p
    ; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5547_clock;
  wire  toggle_5547_reset;
  wire  toggle_5547_valid;
  reg  toggle_5547_valid_reg;
  reg  exu_io_in_bits_r_cf_exceptionVec_2_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  exu_io_in_bits_r_cf_exceptionVec_2_t = exu_io_in_bits_r_cf_exceptionVec_2 ^ exu_io_in_bits_r_cf_exceptionVec_2_p
    ; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5548_clock;
  wire  toggle_5548_reset;
  wire  toggle_5548_valid;
  reg  toggle_5548_valid_reg;
  reg  exu_io_in_bits_r_cf_exceptionVec_12_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  exu_io_in_bits_r_cf_exceptionVec_12_t = exu_io_in_bits_r_cf_exceptionVec_12 ^
    exu_io_in_bits_r_cf_exceptionVec_12_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5549_clock;
  wire  toggle_5549_reset;
  wire  toggle_5549_valid;
  reg  toggle_5549_valid_reg;
  reg  exu_io_in_bits_r_cf_intrVec_1_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  exu_io_in_bits_r_cf_intrVec_1_t = exu_io_in_bits_r_cf_intrVec_1 ^ exu_io_in_bits_r_cf_intrVec_1_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5550_clock;
  wire  toggle_5550_reset;
  wire  toggle_5550_valid;
  reg  toggle_5550_valid_reg;
  reg  exu_io_in_bits_r_cf_intrVec_3_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  exu_io_in_bits_r_cf_intrVec_3_t = exu_io_in_bits_r_cf_intrVec_3 ^ exu_io_in_bits_r_cf_intrVec_3_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5551_clock;
  wire  toggle_5551_reset;
  wire  toggle_5551_valid;
  reg  toggle_5551_valid_reg;
  reg  exu_io_in_bits_r_cf_intrVec_5_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  exu_io_in_bits_r_cf_intrVec_5_t = exu_io_in_bits_r_cf_intrVec_5 ^ exu_io_in_bits_r_cf_intrVec_5_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5552_clock;
  wire  toggle_5552_reset;
  wire  toggle_5552_valid;
  reg  toggle_5552_valid_reg;
  reg  exu_io_in_bits_r_cf_intrVec_7_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  exu_io_in_bits_r_cf_intrVec_7_t = exu_io_in_bits_r_cf_intrVec_7 ^ exu_io_in_bits_r_cf_intrVec_7_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5553_clock;
  wire  toggle_5553_reset;
  wire  toggle_5553_valid;
  reg  toggle_5553_valid_reg;
  reg  exu_io_in_bits_r_cf_intrVec_9_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  exu_io_in_bits_r_cf_intrVec_9_t = exu_io_in_bits_r_cf_intrVec_9 ^ exu_io_in_bits_r_cf_intrVec_9_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5554_clock;
  wire  toggle_5554_reset;
  wire  toggle_5554_valid;
  reg  toggle_5554_valid_reg;
  reg  exu_io_in_bits_r_cf_intrVec_11_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  exu_io_in_bits_r_cf_intrVec_11_t = exu_io_in_bits_r_cf_intrVec_11 ^ exu_io_in_bits_r_cf_intrVec_11_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5555_clock;
  wire  toggle_5555_reset;
  wire  toggle_5555_valid;
  reg  toggle_5555_valid_reg;
  reg [3:0] exu_io_in_bits_r_cf_brIdx_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [3:0] exu_io_in_bits_r_cf_brIdx_t = exu_io_in_bits_r_cf_brIdx ^ exu_io_in_bits_r_cf_brIdx_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5556_clock;
  wire  toggle_5556_reset;
  wire [3:0] toggle_5556_valid;
  reg [3:0] toggle_5556_valid_reg;
  reg  exu_io_in_bits_r_cf_crossBoundaryFault_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  exu_io_in_bits_r_cf_crossBoundaryFault_t = exu_io_in_bits_r_cf_crossBoundaryFault ^
    exu_io_in_bits_r_cf_crossBoundaryFault_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5560_clock;
  wire  toggle_5560_reset;
  wire  toggle_5560_valid;
  reg  toggle_5560_valid_reg;
  reg [2:0] exu_io_in_bits_r_ctrl_fuType_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [2:0] exu_io_in_bits_r_ctrl_fuType_t = exu_io_in_bits_r_ctrl_fuType ^ exu_io_in_bits_r_ctrl_fuType_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5561_clock;
  wire  toggle_5561_reset;
  wire [2:0] toggle_5561_valid;
  reg [2:0] toggle_5561_valid_reg;
  reg [6:0] exu_io_in_bits_r_ctrl_fuOpType_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [6:0] exu_io_in_bits_r_ctrl_fuOpType_t = exu_io_in_bits_r_ctrl_fuOpType ^ exu_io_in_bits_r_ctrl_fuOpType_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5564_clock;
  wire  toggle_5564_reset;
  wire [6:0] toggle_5564_valid;
  reg [6:0] toggle_5564_valid_reg;
  reg  exu_io_in_bits_r_ctrl_rfWen_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  exu_io_in_bits_r_ctrl_rfWen_t = exu_io_in_bits_r_ctrl_rfWen ^ exu_io_in_bits_r_ctrl_rfWen_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5571_clock;
  wire  toggle_5571_reset;
  wire  toggle_5571_valid;
  reg  toggle_5571_valid_reg;
  reg [4:0] exu_io_in_bits_r_ctrl_rfDest_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [4:0] exu_io_in_bits_r_ctrl_rfDest_t = exu_io_in_bits_r_ctrl_rfDest ^ exu_io_in_bits_r_ctrl_rfDest_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5572_clock;
  wire  toggle_5572_reset;
  wire [4:0] toggle_5572_valid;
  reg [4:0] toggle_5572_valid_reg;
  reg  exu_io_in_bits_r_ctrl_isNutCoreTrap_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  exu_io_in_bits_r_ctrl_isNutCoreTrap_t = exu_io_in_bits_r_ctrl_isNutCoreTrap ^
    exu_io_in_bits_r_ctrl_isNutCoreTrap_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5577_clock;
  wire  toggle_5577_reset;
  wire  toggle_5577_valid;
  reg  toggle_5577_valid_reg;
  reg [63:0] exu_io_in_bits_r_data_src1_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [63:0] exu_io_in_bits_r_data_src1_t = exu_io_in_bits_r_data_src1 ^ exu_io_in_bits_r_data_src1_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5578_clock;
  wire  toggle_5578_reset;
  wire [63:0] toggle_5578_valid;
  reg [63:0] toggle_5578_valid_reg;
  reg [63:0] exu_io_in_bits_r_data_src2_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [63:0] exu_io_in_bits_r_data_src2_t = exu_io_in_bits_r_data_src2 ^ exu_io_in_bits_r_data_src2_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5642_clock;
  wire  toggle_5642_reset;
  wire [63:0] toggle_5642_valid;
  reg [63:0] toggle_5642_valid_reg;
  reg [63:0] exu_io_in_bits_r_data_imm_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [63:0] exu_io_in_bits_r_data_imm_t = exu_io_in_bits_r_data_imm ^ exu_io_in_bits_r_data_imm_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5706_clock;
  wire  toggle_5706_reset;
  wire [63:0] toggle_5706_valid;
  reg [63:0] toggle_5706_valid_reg;
  reg  valid_1_p; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  valid_1_t = valid_1 ^ valid_1_p; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  toggle_5770_clock;
  wire  toggle_5770_reset;
  wire  toggle_5770_valid;
  reg  toggle_5770_valid_reg;
  reg [63:0] wbu_io_in_bits_r_decode_cf_instr_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [63:0] wbu_io_in_bits_r_decode_cf_instr_t = wbu_io_in_bits_r_decode_cf_instr ^ wbu_io_in_bits_r_decode_cf_instr_p
    ; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5771_clock;
  wire  toggle_5771_reset;
  wire [63:0] toggle_5771_valid;
  reg [63:0] toggle_5771_valid_reg;
  reg [38:0] wbu_io_in_bits_r_decode_cf_pc_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [38:0] wbu_io_in_bits_r_decode_cf_pc_t = wbu_io_in_bits_r_decode_cf_pc ^ wbu_io_in_bits_r_decode_cf_pc_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5835_clock;
  wire  toggle_5835_reset;
  wire [38:0] toggle_5835_valid;
  reg [38:0] toggle_5835_valid_reg;
  reg [38:0] wbu_io_in_bits_r_decode_cf_redirect_target_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [38:0] wbu_io_in_bits_r_decode_cf_redirect_target_t = wbu_io_in_bits_r_decode_cf_redirect_target ^
    wbu_io_in_bits_r_decode_cf_redirect_target_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5874_clock;
  wire  toggle_5874_reset;
  wire [38:0] toggle_5874_valid;
  reg [38:0] toggle_5874_valid_reg;
  reg  wbu_io_in_bits_r_decode_cf_redirect_valid_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  wbu_io_in_bits_r_decode_cf_redirect_valid_t = wbu_io_in_bits_r_decode_cf_redirect_valid ^
    wbu_io_in_bits_r_decode_cf_redirect_valid_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5913_clock;
  wire  toggle_5913_reset;
  wire  toggle_5913_valid;
  reg  toggle_5913_valid_reg;
  reg [2:0] wbu_io_in_bits_r_decode_ctrl_fuType_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [2:0] wbu_io_in_bits_r_decode_ctrl_fuType_t = wbu_io_in_bits_r_decode_ctrl_fuType ^
    wbu_io_in_bits_r_decode_ctrl_fuType_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5914_clock;
  wire  toggle_5914_reset;
  wire [2:0] toggle_5914_valid;
  reg [2:0] toggle_5914_valid_reg;
  reg  wbu_io_in_bits_r_decode_ctrl_rfWen_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  wbu_io_in_bits_r_decode_ctrl_rfWen_t = wbu_io_in_bits_r_decode_ctrl_rfWen ^ wbu_io_in_bits_r_decode_ctrl_rfWen_p
    ; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5917_clock;
  wire  toggle_5917_reset;
  wire  toggle_5917_valid;
  reg  toggle_5917_valid_reg;
  reg [4:0] wbu_io_in_bits_r_decode_ctrl_rfDest_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [4:0] wbu_io_in_bits_r_decode_ctrl_rfDest_t = wbu_io_in_bits_r_decode_ctrl_rfDest ^
    wbu_io_in_bits_r_decode_ctrl_rfDest_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5918_clock;
  wire  toggle_5918_reset;
  wire [4:0] toggle_5918_valid;
  reg [4:0] toggle_5918_valid_reg;
  reg  wbu_io_in_bits_r_isMMIO_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  wbu_io_in_bits_r_isMMIO_t = wbu_io_in_bits_r_isMMIO ^ wbu_io_in_bits_r_isMMIO_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5923_clock;
  wire  toggle_5923_reset;
  wire  toggle_5923_valid;
  reg  toggle_5923_valid_reg;
  reg [63:0] wbu_io_in_bits_r_commits_0_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [63:0] wbu_io_in_bits_r_commits_0_t = wbu_io_in_bits_r_commits_0 ^ wbu_io_in_bits_r_commits_0_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5924_clock;
  wire  toggle_5924_reset;
  wire [63:0] toggle_5924_valid;
  reg [63:0] toggle_5924_valid_reg;
  reg [63:0] wbu_io_in_bits_r_commits_1_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [63:0] wbu_io_in_bits_r_commits_1_t = wbu_io_in_bits_r_commits_1 ^ wbu_io_in_bits_r_commits_1_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_5988_clock;
  wire  toggle_5988_reset;
  wire [63:0] toggle_5988_valid;
  reg [63:0] toggle_5988_valid_reg;
  reg [63:0] wbu_io_in_bits_r_commits_2_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [63:0] wbu_io_in_bits_r_commits_2_t = wbu_io_in_bits_r_commits_2 ^ wbu_io_in_bits_r_commits_2_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_6052_clock;
  wire  toggle_6052_reset;
  wire [63:0] toggle_6052_valid;
  reg [63:0] toggle_6052_valid_reg;
  reg [63:0] wbu_io_in_bits_r_commits_3_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [63:0] wbu_io_in_bits_r_commits_3_t = wbu_io_in_bits_r_commits_3 ^ wbu_io_in_bits_r_commits_3_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_6116_clock;
  wire  toggle_6116_reset;
  wire [63:0] toggle_6116_valid;
  reg [63:0] toggle_6116_valid_reg;
  reg  wbu_io_in_bits_r_isExit_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  wbu_io_in_bits_r_isExit_t = wbu_io_in_bits_r_isExit ^ wbu_io_in_bits_r_isExit_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_6180_clock;
  wire  toggle_6180_reset;
  wire  toggle_6180_valid;
  reg  toggle_6180_valid_reg;
  ISU isu ( // @[src/main/scala/nutcore/backend/ooo/Backend.scala 679:20]
    .clock(isu_clock),
    .reset(isu_reset),
    .io_in_0_ready(isu_io_in_0_ready),
    .io_in_0_valid(isu_io_in_0_valid),
    .io_in_0_bits_cf_instr(isu_io_in_0_bits_cf_instr),
    .io_in_0_bits_cf_pc(isu_io_in_0_bits_cf_pc),
    .io_in_0_bits_cf_pnpc(isu_io_in_0_bits_cf_pnpc),
    .io_in_0_bits_cf_exceptionVec_1(isu_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(isu_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_exceptionVec_12(isu_io_in_0_bits_cf_exceptionVec_12),
    .io_in_0_bits_cf_intrVec_1(isu_io_in_0_bits_cf_intrVec_1),
    .io_in_0_bits_cf_intrVec_3(isu_io_in_0_bits_cf_intrVec_3),
    .io_in_0_bits_cf_intrVec_5(isu_io_in_0_bits_cf_intrVec_5),
    .io_in_0_bits_cf_intrVec_7(isu_io_in_0_bits_cf_intrVec_7),
    .io_in_0_bits_cf_intrVec_9(isu_io_in_0_bits_cf_intrVec_9),
    .io_in_0_bits_cf_intrVec_11(isu_io_in_0_bits_cf_intrVec_11),
    .io_in_0_bits_cf_brIdx(isu_io_in_0_bits_cf_brIdx),
    .io_in_0_bits_cf_crossBoundaryFault(isu_io_in_0_bits_cf_crossBoundaryFault),
    .io_in_0_bits_ctrl_src1Type(isu_io_in_0_bits_ctrl_src1Type),
    .io_in_0_bits_ctrl_src2Type(isu_io_in_0_bits_ctrl_src2Type),
    .io_in_0_bits_ctrl_fuType(isu_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(isu_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_rfSrc1(isu_io_in_0_bits_ctrl_rfSrc1),
    .io_in_0_bits_ctrl_rfSrc2(isu_io_in_0_bits_ctrl_rfSrc2),
    .io_in_0_bits_ctrl_rfWen(isu_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_rfDest(isu_io_in_0_bits_ctrl_rfDest),
    .io_in_0_bits_ctrl_isNutCoreTrap(isu_io_in_0_bits_ctrl_isNutCoreTrap),
    .io_in_0_bits_data_imm(isu_io_in_0_bits_data_imm),
    .io_out_ready(isu_io_out_ready),
    .io_out_valid(isu_io_out_valid),
    .io_out_bits_cf_instr(isu_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(isu_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(isu_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(isu_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(isu_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_exceptionVec_12(isu_io_out_bits_cf_exceptionVec_12),
    .io_out_bits_cf_intrVec_1(isu_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_3(isu_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_5(isu_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_7(isu_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_9(isu_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_11(isu_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(isu_io_out_bits_cf_brIdx),
    .io_out_bits_cf_crossBoundaryFault(isu_io_out_bits_cf_crossBoundaryFault),
    .io_out_bits_ctrl_fuType(isu_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(isu_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_rfWen(isu_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(isu_io_out_bits_ctrl_rfDest),
    .io_out_bits_ctrl_isNutCoreTrap(isu_io_out_bits_ctrl_isNutCoreTrap),
    .io_out_bits_data_src1(isu_io_out_bits_data_src1),
    .io_out_bits_data_src2(isu_io_out_bits_data_src2),
    .io_out_bits_data_imm(isu_io_out_bits_data_imm),
    .io_wb_rfWen(isu_io_wb_rfWen),
    .io_wb_rfDest(isu_io_wb_rfDest),
    .io_wb_rfData(isu_io_wb_rfData),
    .io_forward_valid(isu_io_forward_valid),
    .io_forward_wb_rfWen(isu_io_forward_wb_rfWen),
    .io_forward_wb_rfDest(isu_io_forward_wb_rfDest),
    .io_forward_wb_rfData(isu_io_forward_wb_rfData),
    .io_forward_fuType(isu_io_forward_fuType),
    .io_flush(isu_io_flush)
  );
  EXU exu ( // @[src/main/scala/nutcore/backend/ooo/Backend.scala 680:20]
    .clock(exu_clock),
    .reset(exu_reset),
    .io__in_ready(exu_io__in_ready),
    .io__in_valid(exu_io__in_valid),
    .io__in_bits_cf_instr(exu_io__in_bits_cf_instr),
    .io__in_bits_cf_pc(exu_io__in_bits_cf_pc),
    .io__in_bits_cf_pnpc(exu_io__in_bits_cf_pnpc),
    .io__in_bits_cf_exceptionVec_1(exu_io__in_bits_cf_exceptionVec_1),
    .io__in_bits_cf_exceptionVec_2(exu_io__in_bits_cf_exceptionVec_2),
    .io__in_bits_cf_exceptionVec_12(exu_io__in_bits_cf_exceptionVec_12),
    .io__in_bits_cf_intrVec_1(exu_io__in_bits_cf_intrVec_1),
    .io__in_bits_cf_intrVec_3(exu_io__in_bits_cf_intrVec_3),
    .io__in_bits_cf_intrVec_5(exu_io__in_bits_cf_intrVec_5),
    .io__in_bits_cf_intrVec_7(exu_io__in_bits_cf_intrVec_7),
    .io__in_bits_cf_intrVec_9(exu_io__in_bits_cf_intrVec_9),
    .io__in_bits_cf_intrVec_11(exu_io__in_bits_cf_intrVec_11),
    .io__in_bits_cf_brIdx(exu_io__in_bits_cf_brIdx),
    .io__in_bits_cf_crossBoundaryFault(exu_io__in_bits_cf_crossBoundaryFault),
    .io__in_bits_ctrl_fuType(exu_io__in_bits_ctrl_fuType),
    .io__in_bits_ctrl_fuOpType(exu_io__in_bits_ctrl_fuOpType),
    .io__in_bits_ctrl_rfWen(exu_io__in_bits_ctrl_rfWen),
    .io__in_bits_ctrl_rfDest(exu_io__in_bits_ctrl_rfDest),
    .io__in_bits_ctrl_isNutCoreTrap(exu_io__in_bits_ctrl_isNutCoreTrap),
    .io__in_bits_data_src1(exu_io__in_bits_data_src1),
    .io__in_bits_data_src2(exu_io__in_bits_data_src2),
    .io__in_bits_data_imm(exu_io__in_bits_data_imm),
    .io__out_ready(exu_io__out_ready),
    .io__out_valid(exu_io__out_valid),
    .io__out_bits_decode_cf_instr(exu_io__out_bits_decode_cf_instr),
    .io__out_bits_decode_cf_pc(exu_io__out_bits_decode_cf_pc),
    .io__out_bits_decode_cf_redirect_target(exu_io__out_bits_decode_cf_redirect_target),
    .io__out_bits_decode_cf_redirect_valid(exu_io__out_bits_decode_cf_redirect_valid),
    .io__out_bits_decode_ctrl_fuType(exu_io__out_bits_decode_ctrl_fuType),
    .io__out_bits_decode_ctrl_rfWen(exu_io__out_bits_decode_ctrl_rfWen),
    .io__out_bits_decode_ctrl_rfDest(exu_io__out_bits_decode_ctrl_rfDest),
    .io__out_bits_isMMIO(exu_io__out_bits_isMMIO),
    .io__out_bits_commits_0(exu_io__out_bits_commits_0),
    .io__out_bits_commits_1(exu_io__out_bits_commits_1),
    .io__out_bits_commits_2(exu_io__out_bits_commits_2),
    .io__out_bits_commits_3(exu_io__out_bits_commits_3),
    .io__out_bits_isExit(exu_io__out_bits_isExit),
    .io__flush(exu_io__flush),
    .io__dmem_req_ready(exu_io__dmem_req_ready),
    .io__dmem_req_valid(exu_io__dmem_req_valid),
    .io__dmem_req_bits_addr(exu_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(exu_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(exu_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(exu_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(exu_io__dmem_req_bits_wdata),
    .io__dmem_resp_valid(exu_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(exu_io__dmem_resp_bits_rdata),
    .io__forward_valid(exu_io__forward_valid),
    .io__forward_wb_rfWen(exu_io__forward_wb_rfWen),
    .io__forward_wb_rfDest(exu_io__forward_wb_rfDest),
    .io__forward_wb_rfData(exu_io__forward_wb_rfData),
    .io__forward_fuType(exu_io__forward_fuType),
    .io__memMMU_imem_priviledgeMode(exu_io__memMMU_imem_priviledgeMode),
    .io__memMMU_dmem_priviledgeMode(exu_io__memMMU_dmem_priviledgeMode),
    .io__memMMU_dmem_status_sum(exu_io__memMMU_dmem_status_sum),
    .io__memMMU_dmem_status_mxr(exu_io__memMMU_dmem_status_mxr),
    .io__memMMU_dmem_loadPF(exu_io__memMMU_dmem_loadPF),
    .io__memMMU_dmem_storePF(exu_io__memMMU_dmem_storePF),
    .io__memMMU_dmem_laf(exu_io__memMMU_dmem_laf),
    .io__memMMU_dmem_saf(exu_io__memMMU_dmem_saf),
    .io__sfence_vma_invalid(exu_io__sfence_vma_invalid),
    .io__wfi_invalid(exu_io__wfi_invalid),
    .lr(exu_lr),
    .io_extra_meip_0(exu_io_extra_meip_0),
    .scInflight(exu_scInflight),
    .REG_valid(exu_REG_valid),
    .REG_pc(exu_REG_pc),
    .REG_isMissPredict(exu_REG_isMissPredict),
    .REG_actualTarget(exu_REG_actualTarget),
    .REG_fuOpType(exu_REG_fuOpType),
    .REG_btbType(exu_REG_btbType),
    .REG_isRVC(exu_REG_isRVC),
    .amoReq(exu_amoReq),
    .lrAddr(exu_lrAddr),
    .paddr(exu_paddr),
    .satp(exu_satp),
    ._T_12_0(exu__T_12_0),
    .scIsSuccess(exu_scIsSuccess),
    .io_extra_mtip(exu_io_extra_mtip),
    .flushICache(exu_flushICache),
    .falseWire(exu_falseWire),
    .vmEnable(exu_vmEnable),
    .flushTLB(exu_flushTLB),
    .intrVecIDU(exu_intrVecIDU),
    .tlbFinish(exu_tlbFinish),
    .ismmio(exu_ismmio),
    ._T_13_1(exu__T_13_1),
    .io_extra_msip(exu_io_extra_msip),
    .io_in_valid(exu_io_in_valid)
  );
  WBU wbu ( // @[src/main/scala/nutcore/backend/ooo/Backend.scala 681:20]
    .clock(wbu_clock),
    .reset(wbu_reset),
    .io__in_valid(wbu_io__in_valid),
    .io__in_bits_decode_cf_instr(wbu_io__in_bits_decode_cf_instr),
    .io__in_bits_decode_cf_pc(wbu_io__in_bits_decode_cf_pc),
    .io__in_bits_decode_cf_redirect_target(wbu_io__in_bits_decode_cf_redirect_target),
    .io__in_bits_decode_cf_redirect_valid(wbu_io__in_bits_decode_cf_redirect_valid),
    .io__in_bits_decode_ctrl_fuType(wbu_io__in_bits_decode_ctrl_fuType),
    .io__in_bits_decode_ctrl_rfWen(wbu_io__in_bits_decode_ctrl_rfWen),
    .io__in_bits_decode_ctrl_rfDest(wbu_io__in_bits_decode_ctrl_rfDest),
    .io__in_bits_isMMIO(wbu_io__in_bits_isMMIO),
    .io__in_bits_commits_0(wbu_io__in_bits_commits_0),
    .io__in_bits_commits_1(wbu_io__in_bits_commits_1),
    .io__in_bits_commits_2(wbu_io__in_bits_commits_2),
    .io__in_bits_commits_3(wbu_io__in_bits_commits_3),
    .io__in_bits_isExit(wbu_io__in_bits_isExit),
    .io__wb_rfWen(wbu_io__wb_rfWen),
    .io__wb_rfDest(wbu_io__wb_rfDest),
    .io__wb_rfData(wbu_io__wb_rfData),
    .io__redirect_target(wbu_io__redirect_target),
    .io__redirect_valid(wbu_io__redirect_valid),
    .falseWire_0(wbu_falseWire_0),
    .io_in_valid(wbu_io_in_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(5404)) toggle_5404 (
    .clock(toggle_5404_clock),
    .reset(toggle_5404_reset),
    .valid(toggle_5404_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(5405)) toggle_5405 (
    .clock(toggle_5405_clock),
    .reset(toggle_5405_reset),
    .valid(toggle_5405_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(5469)) toggle_5469 (
    .clock(toggle_5469_clock),
    .reset(toggle_5469_reset),
    .valid(toggle_5469_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(5508)) toggle_5508 (
    .clock(toggle_5508_clock),
    .reset(toggle_5508_reset),
    .valid(toggle_5508_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(5547)) toggle_5547 (
    .clock(toggle_5547_clock),
    .reset(toggle_5547_reset),
    .valid(toggle_5547_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(5548)) toggle_5548 (
    .clock(toggle_5548_clock),
    .reset(toggle_5548_reset),
    .valid(toggle_5548_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(5549)) toggle_5549 (
    .clock(toggle_5549_clock),
    .reset(toggle_5549_reset),
    .valid(toggle_5549_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(5550)) toggle_5550 (
    .clock(toggle_5550_clock),
    .reset(toggle_5550_reset),
    .valid(toggle_5550_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(5551)) toggle_5551 (
    .clock(toggle_5551_clock),
    .reset(toggle_5551_reset),
    .valid(toggle_5551_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(5552)) toggle_5552 (
    .clock(toggle_5552_clock),
    .reset(toggle_5552_reset),
    .valid(toggle_5552_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(5553)) toggle_5553 (
    .clock(toggle_5553_clock),
    .reset(toggle_5553_reset),
    .valid(toggle_5553_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(5554)) toggle_5554 (
    .clock(toggle_5554_clock),
    .reset(toggle_5554_reset),
    .valid(toggle_5554_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(5555)) toggle_5555 (
    .clock(toggle_5555_clock),
    .reset(toggle_5555_reset),
    .valid(toggle_5555_valid)
  );
  GEN_w4_toggle #(.COVER_INDEX(5556)) toggle_5556 (
    .clock(toggle_5556_clock),
    .reset(toggle_5556_reset),
    .valid(toggle_5556_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(5560)) toggle_5560 (
    .clock(toggle_5560_clock),
    .reset(toggle_5560_reset),
    .valid(toggle_5560_valid)
  );
  GEN_w3_toggle #(.COVER_INDEX(5561)) toggle_5561 (
    .clock(toggle_5561_clock),
    .reset(toggle_5561_reset),
    .valid(toggle_5561_valid)
  );
  GEN_w7_toggle #(.COVER_INDEX(5564)) toggle_5564 (
    .clock(toggle_5564_clock),
    .reset(toggle_5564_reset),
    .valid(toggle_5564_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(5571)) toggle_5571 (
    .clock(toggle_5571_clock),
    .reset(toggle_5571_reset),
    .valid(toggle_5571_valid)
  );
  GEN_w5_toggle #(.COVER_INDEX(5572)) toggle_5572 (
    .clock(toggle_5572_clock),
    .reset(toggle_5572_reset),
    .valid(toggle_5572_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(5577)) toggle_5577 (
    .clock(toggle_5577_clock),
    .reset(toggle_5577_reset),
    .valid(toggle_5577_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(5578)) toggle_5578 (
    .clock(toggle_5578_clock),
    .reset(toggle_5578_reset),
    .valid(toggle_5578_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(5642)) toggle_5642 (
    .clock(toggle_5642_clock),
    .reset(toggle_5642_reset),
    .valid(toggle_5642_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(5706)) toggle_5706 (
    .clock(toggle_5706_clock),
    .reset(toggle_5706_reset),
    .valid(toggle_5706_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(5770)) toggle_5770 (
    .clock(toggle_5770_clock),
    .reset(toggle_5770_reset),
    .valid(toggle_5770_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(5771)) toggle_5771 (
    .clock(toggle_5771_clock),
    .reset(toggle_5771_reset),
    .valid(toggle_5771_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(5835)) toggle_5835 (
    .clock(toggle_5835_clock),
    .reset(toggle_5835_reset),
    .valid(toggle_5835_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(5874)) toggle_5874 (
    .clock(toggle_5874_clock),
    .reset(toggle_5874_reset),
    .valid(toggle_5874_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(5913)) toggle_5913 (
    .clock(toggle_5913_clock),
    .reset(toggle_5913_reset),
    .valid(toggle_5913_valid)
  );
  GEN_w3_toggle #(.COVER_INDEX(5914)) toggle_5914 (
    .clock(toggle_5914_clock),
    .reset(toggle_5914_reset),
    .valid(toggle_5914_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(5917)) toggle_5917 (
    .clock(toggle_5917_clock),
    .reset(toggle_5917_reset),
    .valid(toggle_5917_valid)
  );
  GEN_w5_toggle #(.COVER_INDEX(5918)) toggle_5918 (
    .clock(toggle_5918_clock),
    .reset(toggle_5918_reset),
    .valid(toggle_5918_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(5923)) toggle_5923 (
    .clock(toggle_5923_clock),
    .reset(toggle_5923_reset),
    .valid(toggle_5923_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(5924)) toggle_5924 (
    .clock(toggle_5924_clock),
    .reset(toggle_5924_reset),
    .valid(toggle_5924_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(5988)) toggle_5988 (
    .clock(toggle_5988_clock),
    .reset(toggle_5988_reset),
    .valid(toggle_5988_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(6052)) toggle_6052 (
    .clock(toggle_6052_clock),
    .reset(toggle_6052_reset),
    .valid(toggle_6052_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(6116)) toggle_6116 (
    .clock(toggle_6116_clock),
    .reset(toggle_6116_reset),
    .valid(toggle_6116_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(6180)) toggle_6180 (
    .clock(toggle_6180_clock),
    .reset(toggle_6180_reset),
    .valid(toggle_6180_valid)
  );
  assign io_in_0_ready = isu_io_in_0_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign io_dmem_req_valid = exu_io__dmem_req_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign io_dmem_req_bits_addr = exu_io__dmem_req_bits_addr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign io_dmem_req_bits_size = exu_io__dmem_req_bits_size; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign io_dmem_req_bits_cmd = exu_io__dmem_req_bits_cmd; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign io_dmem_req_bits_wmask = exu_io__dmem_req_bits_wmask; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign io_dmem_req_bits_wdata = exu_io__dmem_req_bits_wdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign io_memMMU_imem_priviledgeMode = exu_io__memMMU_imem_priviledgeMode; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 698:18]
  assign io_memMMU_dmem_priviledgeMode = exu_io__memMMU_dmem_priviledgeMode; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign io_memMMU_dmem_status_sum = exu_io__memMMU_dmem_status_sum; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign io_memMMU_dmem_status_mxr = exu_io__memMMU_dmem_status_mxr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign io_sfence_vma_invalid = exu_io__sfence_vma_invalid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 692:25]
  assign io_wfi_invalid = exu_io__wfi_invalid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 693:18]
  assign io_redirect_target = wbu_io__redirect_target; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 694:15]
  assign io_redirect_valid = wbu_io__redirect_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 694:15]
  assign lr = exu_lr;
  assign scInflight = exu_scInflight;
  assign REG_valid = exu_REG_valid;
  assign REG_pc = exu_REG_pc;
  assign REG_isMissPredict = exu_REG_isMissPredict;
  assign REG_actualTarget = exu_REG_actualTarget;
  assign REG_fuOpType = exu_REG_fuOpType;
  assign REG_btbType = exu_REG_btbType;
  assign REG_isRVC = exu_REG_isRVC;
  assign amoReq = exu_amoReq;
  assign lrAddr = exu_lrAddr;
  assign satp = exu_satp;
  assign flushICache = exu_flushICache;
  assign flushTLB = exu_flushTLB;
  assign intrVecIDU = exu_intrVecIDU;
  assign isu_clock = clock;
  assign isu_reset = reset;
  assign isu_io_in_0_valid = io_in_0_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_instr = io_in_0_bits_cf_instr; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_pc = io_in_0_bits_cf_pc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_pnpc = io_in_0_bits_cf_pnpc; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_exceptionVec_1 = io_in_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_exceptionVec_2 = io_in_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_exceptionVec_12 = io_in_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_intrVec_1 = io_in_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_intrVec_3 = io_in_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_intrVec_5 = io_in_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_intrVec_7 = io_in_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_intrVec_9 = io_in_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_intrVec_11 = io_in_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_brIdx = io_in_0_bits_cf_brIdx; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_cf_crossBoundaryFault = io_in_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_src1Type = io_in_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_src2Type = io_in_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_fuType = io_in_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_fuOpType = io_in_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_rfSrc1 = io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_rfSrc2 = io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_rfWen = io_in_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_rfDest = io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_ctrl_isNutCoreTrap = io_in_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_in_0_bits_data_imm = io_in_0_bits_data_imm; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 686:13]
  assign isu_io_out_ready = exu_io__in_ready; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign isu_io_wb_rfWen = wbu_io__wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 691:13]
  assign isu_io_wb_rfDest = wbu_io__wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 691:13]
  assign isu_io_wb_rfData = wbu_io__wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 691:13]
  assign isu_io_forward_valid = exu_io__forward_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign isu_io_forward_wb_rfWen = exu_io__forward_wb_rfWen; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign isu_io_forward_wb_rfDest = exu_io__forward_wb_rfDest; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign isu_io_forward_wb_rfData = exu_io__forward_wb_rfData; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign isu_io_forward_fuType = exu_io__forward_fuType; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 696:18]
  assign isu_io_flush = io_flush[0]; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 688:27]
  assign exu_clock = clock;
  assign exu_reset = reset;
  assign exu_io__in_valid = valid; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign exu_io__in_bits_cf_instr = exu_io_in_bits_r_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_pc = exu_io_in_bits_r_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_pnpc = exu_io_in_bits_r_cf_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_1 = exu_io_in_bits_r_cf_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_2 = exu_io_in_bits_r_cf_exceptionVec_2; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_12 = exu_io_in_bits_r_cf_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_1 = exu_io_in_bits_r_cf_intrVec_1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_3 = exu_io_in_bits_r_cf_intrVec_3; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_5 = exu_io_in_bits_r_cf_intrVec_5; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_7 = exu_io_in_bits_r_cf_intrVec_7; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_9 = exu_io_in_bits_r_cf_intrVec_9; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_11 = exu_io_in_bits_r_cf_intrVec_11; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_brIdx = exu_io_in_bits_r_cf_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_crossBoundaryFault = exu_io_in_bits_r_cf_crossBoundaryFault; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_fuType = exu_io_in_bits_r_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_fuOpType = exu_io_in_bits_r_ctrl_fuOpType; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_rfWen = exu_io_in_bits_r_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_rfDest = exu_io_in_bits_r_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_isNutCoreTrap = exu_io_in_bits_r_ctrl_isNutCoreTrap; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_data_src1 = exu_io_in_bits_r_data_src1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_data_src2 = exu_io_in_bits_r_data_src2; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__in_bits_data_imm = exu_io_in_bits_r_data_imm; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign exu_io__out_ready = 1'h1; // @[src/main/scala/utils/Pipeline.scala 29:16]
  assign exu_io__flush = io_flush[1]; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 689:27]
  assign exu_io__dmem_req_ready = io_dmem_req_ready; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign exu_io__dmem_resp_valid = io_dmem_resp_valid; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign exu_io__dmem_resp_bits_rdata = io_dmem_resp_bits_rdata; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 700:11]
  assign exu_io__memMMU_dmem_loadPF = io_memMMU_dmem_loadPF; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign exu_io__memMMU_dmem_storePF = io_memMMU_dmem_storePF; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign exu_io__memMMU_dmem_laf = io_memMMU_dmem_laf; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign exu_io__memMMU_dmem_saf = io_memMMU_dmem_saf; // @[src/main/scala/nutcore/backend/ooo/Backend.scala 699:18]
  assign exu_io_extra_meip_0 = io_extra_meip_0;
  assign exu_paddr = paddr;
  assign exu__T_12_0 = _T_12;
  assign exu_scIsSuccess = scIsSuccess;
  assign exu_io_extra_mtip = io_extra_mtip;
  assign exu_falseWire = wbu_falseWire_0;
  assign exu_vmEnable = vmEnable;
  assign exu_tlbFinish = tlbFinish;
  assign exu_ismmio = ismmio;
  assign exu__T_13_1 = _T_13_0;
  assign exu_io_extra_msip = io_extra_msip;
  assign exu_io_in_valid = wbu_io_in_valid;
  assign wbu_clock = clock;
  assign wbu_reset = reset;
  assign wbu_io__in_valid = valid_1; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign wbu_io__in_bits_decode_cf_instr = wbu_io_in_bits_r_decode_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_pc = wbu_io_in_bits_r_decode_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_redirect_target = wbu_io_in_bits_r_decode_cf_redirect_target; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_redirect_valid = wbu_io_in_bits_r_decode_cf_redirect_valid; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_fuType = wbu_io_in_bits_r_decode_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_rfWen = wbu_io_in_bits_r_decode_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_rfDest = wbu_io_in_bits_r_decode_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_isMMIO = wbu_io_in_bits_r_isMMIO; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_0 = wbu_io_in_bits_r_commits_0; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_1 = wbu_io_in_bits_r_commits_1; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_2 = wbu_io_in_bits_r_commits_2; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_3 = wbu_io_in_bits_r_commits_3; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign wbu_io__in_bits_isExit = wbu_io_in_bits_r_isExit; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign toggle_5404_clock = clock;
  assign toggle_5404_reset = reset;
  assign toggle_5404_valid = valid ^ toggle_5404_valid_reg;
  assign toggle_5405_clock = clock;
  assign toggle_5405_reset = reset;
  assign toggle_5405_valid = exu_io_in_bits_r_cf_instr ^ toggle_5405_valid_reg;
  assign toggle_5469_clock = clock;
  assign toggle_5469_reset = reset;
  assign toggle_5469_valid = exu_io_in_bits_r_cf_pc ^ toggle_5469_valid_reg;
  assign toggle_5508_clock = clock;
  assign toggle_5508_reset = reset;
  assign toggle_5508_valid = exu_io_in_bits_r_cf_pnpc ^ toggle_5508_valid_reg;
  assign toggle_5547_clock = clock;
  assign toggle_5547_reset = reset;
  assign toggle_5547_valid = exu_io_in_bits_r_cf_exceptionVec_1 ^ toggle_5547_valid_reg;
  assign toggle_5548_clock = clock;
  assign toggle_5548_reset = reset;
  assign toggle_5548_valid = exu_io_in_bits_r_cf_exceptionVec_2 ^ toggle_5548_valid_reg;
  assign toggle_5549_clock = clock;
  assign toggle_5549_reset = reset;
  assign toggle_5549_valid = exu_io_in_bits_r_cf_exceptionVec_12 ^ toggle_5549_valid_reg;
  assign toggle_5550_clock = clock;
  assign toggle_5550_reset = reset;
  assign toggle_5550_valid = exu_io_in_bits_r_cf_intrVec_1 ^ toggle_5550_valid_reg;
  assign toggle_5551_clock = clock;
  assign toggle_5551_reset = reset;
  assign toggle_5551_valid = exu_io_in_bits_r_cf_intrVec_3 ^ toggle_5551_valid_reg;
  assign toggle_5552_clock = clock;
  assign toggle_5552_reset = reset;
  assign toggle_5552_valid = exu_io_in_bits_r_cf_intrVec_5 ^ toggle_5552_valid_reg;
  assign toggle_5553_clock = clock;
  assign toggle_5553_reset = reset;
  assign toggle_5553_valid = exu_io_in_bits_r_cf_intrVec_7 ^ toggle_5553_valid_reg;
  assign toggle_5554_clock = clock;
  assign toggle_5554_reset = reset;
  assign toggle_5554_valid = exu_io_in_bits_r_cf_intrVec_9 ^ toggle_5554_valid_reg;
  assign toggle_5555_clock = clock;
  assign toggle_5555_reset = reset;
  assign toggle_5555_valid = exu_io_in_bits_r_cf_intrVec_11 ^ toggle_5555_valid_reg;
  assign toggle_5556_clock = clock;
  assign toggle_5556_reset = reset;
  assign toggle_5556_valid = exu_io_in_bits_r_cf_brIdx ^ toggle_5556_valid_reg;
  assign toggle_5560_clock = clock;
  assign toggle_5560_reset = reset;
  assign toggle_5560_valid = exu_io_in_bits_r_cf_crossBoundaryFault ^ toggle_5560_valid_reg;
  assign toggle_5561_clock = clock;
  assign toggle_5561_reset = reset;
  assign toggle_5561_valid = exu_io_in_bits_r_ctrl_fuType ^ toggle_5561_valid_reg;
  assign toggle_5564_clock = clock;
  assign toggle_5564_reset = reset;
  assign toggle_5564_valid = exu_io_in_bits_r_ctrl_fuOpType ^ toggle_5564_valid_reg;
  assign toggle_5571_clock = clock;
  assign toggle_5571_reset = reset;
  assign toggle_5571_valid = exu_io_in_bits_r_ctrl_rfWen ^ toggle_5571_valid_reg;
  assign toggle_5572_clock = clock;
  assign toggle_5572_reset = reset;
  assign toggle_5572_valid = exu_io_in_bits_r_ctrl_rfDest ^ toggle_5572_valid_reg;
  assign toggle_5577_clock = clock;
  assign toggle_5577_reset = reset;
  assign toggle_5577_valid = exu_io_in_bits_r_ctrl_isNutCoreTrap ^ toggle_5577_valid_reg;
  assign toggle_5578_clock = clock;
  assign toggle_5578_reset = reset;
  assign toggle_5578_valid = exu_io_in_bits_r_data_src1 ^ toggle_5578_valid_reg;
  assign toggle_5642_clock = clock;
  assign toggle_5642_reset = reset;
  assign toggle_5642_valid = exu_io_in_bits_r_data_src2 ^ toggle_5642_valid_reg;
  assign toggle_5706_clock = clock;
  assign toggle_5706_reset = reset;
  assign toggle_5706_valid = exu_io_in_bits_r_data_imm ^ toggle_5706_valid_reg;
  assign toggle_5770_clock = clock;
  assign toggle_5770_reset = reset;
  assign toggle_5770_valid = valid_1 ^ toggle_5770_valid_reg;
  assign toggle_5771_clock = clock;
  assign toggle_5771_reset = reset;
  assign toggle_5771_valid = wbu_io_in_bits_r_decode_cf_instr ^ toggle_5771_valid_reg;
  assign toggle_5835_clock = clock;
  assign toggle_5835_reset = reset;
  assign toggle_5835_valid = wbu_io_in_bits_r_decode_cf_pc ^ toggle_5835_valid_reg;
  assign toggle_5874_clock = clock;
  assign toggle_5874_reset = reset;
  assign toggle_5874_valid = wbu_io_in_bits_r_decode_cf_redirect_target ^ toggle_5874_valid_reg;
  assign toggle_5913_clock = clock;
  assign toggle_5913_reset = reset;
  assign toggle_5913_valid = wbu_io_in_bits_r_decode_cf_redirect_valid ^ toggle_5913_valid_reg;
  assign toggle_5914_clock = clock;
  assign toggle_5914_reset = reset;
  assign toggle_5914_valid = wbu_io_in_bits_r_decode_ctrl_fuType ^ toggle_5914_valid_reg;
  assign toggle_5917_clock = clock;
  assign toggle_5917_reset = reset;
  assign toggle_5917_valid = wbu_io_in_bits_r_decode_ctrl_rfWen ^ toggle_5917_valid_reg;
  assign toggle_5918_clock = clock;
  assign toggle_5918_reset = reset;
  assign toggle_5918_valid = wbu_io_in_bits_r_decode_ctrl_rfDest ^ toggle_5918_valid_reg;
  assign toggle_5923_clock = clock;
  assign toggle_5923_reset = reset;
  assign toggle_5923_valid = wbu_io_in_bits_r_isMMIO ^ toggle_5923_valid_reg;
  assign toggle_5924_clock = clock;
  assign toggle_5924_reset = reset;
  assign toggle_5924_valid = wbu_io_in_bits_r_commits_0 ^ toggle_5924_valid_reg;
  assign toggle_5988_clock = clock;
  assign toggle_5988_reset = reset;
  assign toggle_5988_valid = wbu_io_in_bits_r_commits_1 ^ toggle_5988_valid_reg;
  assign toggle_6052_clock = clock;
  assign toggle_6052_reset = reset;
  assign toggle_6052_valid = wbu_io_in_bits_r_commits_2 ^ toggle_6052_valid_reg;
  assign toggle_6116_clock = clock;
  assign toggle_6116_reset = reset;
  assign toggle_6116_valid = wbu_io_in_bits_r_commits_3 ^ toggle_6116_valid_reg;
  assign toggle_6180_clock = clock;
  assign toggle_6180_reset = reset;
  assign toggle_6180_valid = wbu_io_in_bits_r_isExit ^ toggle_6180_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else if (io_flush[0]) begin // @[src/main/scala/utils/Pipeline.scala 27:20]
      valid <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 27:28]
    end else begin
      valid <= _GEN_1;
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_instr <= isu_io_out_bits_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_pc <= isu_io_out_bits_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_pnpc <= isu_io_out_bits_cf_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_exceptionVec_1 <= isu_io_out_bits_cf_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_exceptionVec_2 <= isu_io_out_bits_cf_exceptionVec_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_exceptionVec_12 <= isu_io_out_bits_cf_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_1 <= isu_io_out_bits_cf_intrVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_3 <= isu_io_out_bits_cf_intrVec_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_5 <= isu_io_out_bits_cf_intrVec_5; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_7 <= isu_io_out_bits_cf_intrVec_7; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_9 <= isu_io_out_bits_cf_intrVec_9; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_intrVec_11 <= isu_io_out_bits_cf_intrVec_11; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_brIdx <= isu_io_out_bits_cf_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_cf_crossBoundaryFault <= isu_io_out_bits_cf_crossBoundaryFault; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_fuType <= isu_io_out_bits_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_fuOpType <= isu_io_out_bits_ctrl_fuOpType; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_rfWen <= isu_io_out_bits_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_rfDest <= isu_io_out_bits_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_ctrl_isNutCoreTrap <= isu_io_out_bits_ctrl_isNutCoreTrap; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_data_src1 <= isu_io_out_bits_data_src1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_data_src2 <= isu_io_out_bits_data_src2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_2) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      exu_io_in_bits_r_data_imm <= isu_io_out_bits_data_imm; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid_1 <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else if (io_flush[1]) begin // @[src/main/scala/utils/Pipeline.scala 27:20]
      valid_1 <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 27:28]
    end else begin
      valid_1 <= _T_4;
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_cf_instr <= exu_io__out_bits_decode_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_cf_pc <= exu_io__out_bits_decode_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_cf_redirect_target <= exu_io__out_bits_decode_cf_redirect_target; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_cf_redirect_valid <= exu_io__out_bits_decode_cf_redirect_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_ctrl_fuType <= exu_io__out_bits_decode_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_ctrl_rfWen <= exu_io__out_bits_decode_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_decode_ctrl_rfDest <= exu_io__out_bits_decode_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_isMMIO <= exu_io__out_bits_isMMIO; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_commits_0 <= exu_io__out_bits_commits_0; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_commits_1 <= exu_io__out_bits_commits_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_commits_2 <= exu_io__out_bits_commits_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_commits_3 <= exu_io__out_bits_commits_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_4) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      wbu_io_in_bits_r_isExit <= exu_io__out_bits_isExit; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    valid_p <= valid; // @[src/main/scala/utils/Pipeline.scala 24:24]
    toggle_5404_valid_reg <= valid;
    exu_io_in_bits_r_cf_instr_p <= exu_io_in_bits_r_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5405_valid_reg <= exu_io_in_bits_r_cf_instr;
    exu_io_in_bits_r_cf_pc_p <= exu_io_in_bits_r_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5469_valid_reg <= exu_io_in_bits_r_cf_pc;
    exu_io_in_bits_r_cf_pnpc_p <= exu_io_in_bits_r_cf_pnpc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5508_valid_reg <= exu_io_in_bits_r_cf_pnpc;
    exu_io_in_bits_r_cf_exceptionVec_1_p <= exu_io_in_bits_r_cf_exceptionVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5547_valid_reg <= exu_io_in_bits_r_cf_exceptionVec_1;
    exu_io_in_bits_r_cf_exceptionVec_2_p <= exu_io_in_bits_r_cf_exceptionVec_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5548_valid_reg <= exu_io_in_bits_r_cf_exceptionVec_2;
    exu_io_in_bits_r_cf_exceptionVec_12_p <= exu_io_in_bits_r_cf_exceptionVec_12; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5549_valid_reg <= exu_io_in_bits_r_cf_exceptionVec_12;
    exu_io_in_bits_r_cf_intrVec_1_p <= exu_io_in_bits_r_cf_intrVec_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5550_valid_reg <= exu_io_in_bits_r_cf_intrVec_1;
    exu_io_in_bits_r_cf_intrVec_3_p <= exu_io_in_bits_r_cf_intrVec_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5551_valid_reg <= exu_io_in_bits_r_cf_intrVec_3;
    exu_io_in_bits_r_cf_intrVec_5_p <= exu_io_in_bits_r_cf_intrVec_5; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5552_valid_reg <= exu_io_in_bits_r_cf_intrVec_5;
    exu_io_in_bits_r_cf_intrVec_7_p <= exu_io_in_bits_r_cf_intrVec_7; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5553_valid_reg <= exu_io_in_bits_r_cf_intrVec_7;
    exu_io_in_bits_r_cf_intrVec_9_p <= exu_io_in_bits_r_cf_intrVec_9; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5554_valid_reg <= exu_io_in_bits_r_cf_intrVec_9;
    exu_io_in_bits_r_cf_intrVec_11_p <= exu_io_in_bits_r_cf_intrVec_11; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5555_valid_reg <= exu_io_in_bits_r_cf_intrVec_11;
    exu_io_in_bits_r_cf_brIdx_p <= exu_io_in_bits_r_cf_brIdx; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5556_valid_reg <= exu_io_in_bits_r_cf_brIdx;
    exu_io_in_bits_r_cf_crossBoundaryFault_p <= exu_io_in_bits_r_cf_crossBoundaryFault; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5560_valid_reg <= exu_io_in_bits_r_cf_crossBoundaryFault;
    exu_io_in_bits_r_ctrl_fuType_p <= exu_io_in_bits_r_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5561_valid_reg <= exu_io_in_bits_r_ctrl_fuType;
    exu_io_in_bits_r_ctrl_fuOpType_p <= exu_io_in_bits_r_ctrl_fuOpType; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5564_valid_reg <= exu_io_in_bits_r_ctrl_fuOpType;
    exu_io_in_bits_r_ctrl_rfWen_p <= exu_io_in_bits_r_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5571_valid_reg <= exu_io_in_bits_r_ctrl_rfWen;
    exu_io_in_bits_r_ctrl_rfDest_p <= exu_io_in_bits_r_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5572_valid_reg <= exu_io_in_bits_r_ctrl_rfDest;
    exu_io_in_bits_r_ctrl_isNutCoreTrap_p <= exu_io_in_bits_r_ctrl_isNutCoreTrap; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5577_valid_reg <= exu_io_in_bits_r_ctrl_isNutCoreTrap;
    exu_io_in_bits_r_data_src1_p <= exu_io_in_bits_r_data_src1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5578_valid_reg <= exu_io_in_bits_r_data_src1;
    exu_io_in_bits_r_data_src2_p <= exu_io_in_bits_r_data_src2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5642_valid_reg <= exu_io_in_bits_r_data_src2;
    exu_io_in_bits_r_data_imm_p <= exu_io_in_bits_r_data_imm; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5706_valid_reg <= exu_io_in_bits_r_data_imm;
    valid_1_p <= valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24]
    toggle_5770_valid_reg <= valid_1;
    wbu_io_in_bits_r_decode_cf_instr_p <= wbu_io_in_bits_r_decode_cf_instr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5771_valid_reg <= wbu_io_in_bits_r_decode_cf_instr;
    wbu_io_in_bits_r_decode_cf_pc_p <= wbu_io_in_bits_r_decode_cf_pc; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5835_valid_reg <= wbu_io_in_bits_r_decode_cf_pc;
    wbu_io_in_bits_r_decode_cf_redirect_target_p <= wbu_io_in_bits_r_decode_cf_redirect_target; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5874_valid_reg <= wbu_io_in_bits_r_decode_cf_redirect_target;
    wbu_io_in_bits_r_decode_cf_redirect_valid_p <= wbu_io_in_bits_r_decode_cf_redirect_valid; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5913_valid_reg <= wbu_io_in_bits_r_decode_cf_redirect_valid;
    wbu_io_in_bits_r_decode_ctrl_fuType_p <= wbu_io_in_bits_r_decode_ctrl_fuType; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5914_valid_reg <= wbu_io_in_bits_r_decode_ctrl_fuType;
    wbu_io_in_bits_r_decode_ctrl_rfWen_p <= wbu_io_in_bits_r_decode_ctrl_rfWen; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5917_valid_reg <= wbu_io_in_bits_r_decode_ctrl_rfWen;
    wbu_io_in_bits_r_decode_ctrl_rfDest_p <= wbu_io_in_bits_r_decode_ctrl_rfDest; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5918_valid_reg <= wbu_io_in_bits_r_decode_ctrl_rfDest;
    wbu_io_in_bits_r_isMMIO_p <= wbu_io_in_bits_r_isMMIO; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5923_valid_reg <= wbu_io_in_bits_r_isMMIO;
    wbu_io_in_bits_r_commits_0_p <= wbu_io_in_bits_r_commits_0; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5924_valid_reg <= wbu_io_in_bits_r_commits_0;
    wbu_io_in_bits_r_commits_1_p <= wbu_io_in_bits_r_commits_1; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_5988_valid_reg <= wbu_io_in_bits_r_commits_1;
    wbu_io_in_bits_r_commits_2_p <= wbu_io_in_bits_r_commits_2; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_6052_valid_reg <= wbu_io_in_bits_r_commits_2;
    wbu_io_in_bits_r_commits_3_p <= wbu_io_in_bits_r_commits_3; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_6116_valid_reg <= wbu_io_in_bits_r_commits_3;
    wbu_io_in_bits_r_isExit_p <= wbu_io_in_bits_r_isExit; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_6180_valid_reg <= wbu_io_in_bits_r_isExit;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  exu_io_in_bits_r_cf_instr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  exu_io_in_bits_r_cf_pc = _RAND_2[38:0];
  _RAND_3 = {2{`RANDOM}};
  exu_io_in_bits_r_cf_pnpc = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_exceptionVec_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_exceptionVec_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_exceptionVec_12 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_5 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_7 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_9 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_11 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_brIdx = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_crossBoundaryFault = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_fuType = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_fuOpType = _RAND_16[6:0];
  _RAND_17 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_rfWen = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_rfDest = _RAND_18[4:0];
  _RAND_19 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_isNutCoreTrap = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  exu_io_in_bits_r_data_src1 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  exu_io_in_bits_r_data_src2 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  exu_io_in_bits_r_data_imm = _RAND_22[63:0];
  _RAND_23 = {1{`RANDOM}};
  valid_1 = _RAND_23[0:0];
  _RAND_24 = {2{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_instr = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_pc = _RAND_25[38:0];
  _RAND_26 = {2{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_redirect_target = _RAND_26[38:0];
  _RAND_27 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_redirect_valid = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_ctrl_fuType = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_ctrl_rfWen = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_ctrl_rfDest = _RAND_30[4:0];
  _RAND_31 = {1{`RANDOM}};
  wbu_io_in_bits_r_isMMIO = _RAND_31[0:0];
  _RAND_32 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_0 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_1 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_2 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_3 = _RAND_35[63:0];
  _RAND_36 = {1{`RANDOM}};
  wbu_io_in_bits_r_isExit = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  valid_p = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  toggle_5404_valid_reg = _RAND_38[0:0];
  _RAND_39 = {2{`RANDOM}};
  exu_io_in_bits_r_cf_instr_p = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  toggle_5405_valid_reg = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  exu_io_in_bits_r_cf_pc_p = _RAND_41[38:0];
  _RAND_42 = {2{`RANDOM}};
  toggle_5469_valid_reg = _RAND_42[38:0];
  _RAND_43 = {2{`RANDOM}};
  exu_io_in_bits_r_cf_pnpc_p = _RAND_43[38:0];
  _RAND_44 = {2{`RANDOM}};
  toggle_5508_valid_reg = _RAND_44[38:0];
  _RAND_45 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_exceptionVec_1_p = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  toggle_5547_valid_reg = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_exceptionVec_2_p = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  toggle_5548_valid_reg = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_exceptionVec_12_p = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  toggle_5549_valid_reg = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_1_p = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  toggle_5550_valid_reg = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_3_p = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  toggle_5551_valid_reg = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_5_p = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  toggle_5552_valid_reg = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_7_p = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  toggle_5553_valid_reg = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_9_p = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  toggle_5554_valid_reg = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_intrVec_11_p = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  toggle_5555_valid_reg = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_brIdx_p = _RAND_63[3:0];
  _RAND_64 = {1{`RANDOM}};
  toggle_5556_valid_reg = _RAND_64[3:0];
  _RAND_65 = {1{`RANDOM}};
  exu_io_in_bits_r_cf_crossBoundaryFault_p = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  toggle_5560_valid_reg = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_fuType_p = _RAND_67[2:0];
  _RAND_68 = {1{`RANDOM}};
  toggle_5561_valid_reg = _RAND_68[2:0];
  _RAND_69 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_fuOpType_p = _RAND_69[6:0];
  _RAND_70 = {1{`RANDOM}};
  toggle_5564_valid_reg = _RAND_70[6:0];
  _RAND_71 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_rfWen_p = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  toggle_5571_valid_reg = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_rfDest_p = _RAND_73[4:0];
  _RAND_74 = {1{`RANDOM}};
  toggle_5572_valid_reg = _RAND_74[4:0];
  _RAND_75 = {1{`RANDOM}};
  exu_io_in_bits_r_ctrl_isNutCoreTrap_p = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  toggle_5577_valid_reg = _RAND_76[0:0];
  _RAND_77 = {2{`RANDOM}};
  exu_io_in_bits_r_data_src1_p = _RAND_77[63:0];
  _RAND_78 = {2{`RANDOM}};
  toggle_5578_valid_reg = _RAND_78[63:0];
  _RAND_79 = {2{`RANDOM}};
  exu_io_in_bits_r_data_src2_p = _RAND_79[63:0];
  _RAND_80 = {2{`RANDOM}};
  toggle_5642_valid_reg = _RAND_80[63:0];
  _RAND_81 = {2{`RANDOM}};
  exu_io_in_bits_r_data_imm_p = _RAND_81[63:0];
  _RAND_82 = {2{`RANDOM}};
  toggle_5706_valid_reg = _RAND_82[63:0];
  _RAND_83 = {1{`RANDOM}};
  valid_1_p = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  toggle_5770_valid_reg = _RAND_84[0:0];
  _RAND_85 = {2{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_instr_p = _RAND_85[63:0];
  _RAND_86 = {2{`RANDOM}};
  toggle_5771_valid_reg = _RAND_86[63:0];
  _RAND_87 = {2{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_pc_p = _RAND_87[38:0];
  _RAND_88 = {2{`RANDOM}};
  toggle_5835_valid_reg = _RAND_88[38:0];
  _RAND_89 = {2{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_redirect_target_p = _RAND_89[38:0];
  _RAND_90 = {2{`RANDOM}};
  toggle_5874_valid_reg = _RAND_90[38:0];
  _RAND_91 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_cf_redirect_valid_p = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  toggle_5913_valid_reg = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_ctrl_fuType_p = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  toggle_5914_valid_reg = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_ctrl_rfWen_p = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  toggle_5917_valid_reg = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  wbu_io_in_bits_r_decode_ctrl_rfDest_p = _RAND_97[4:0];
  _RAND_98 = {1{`RANDOM}};
  toggle_5918_valid_reg = _RAND_98[4:0];
  _RAND_99 = {1{`RANDOM}};
  wbu_io_in_bits_r_isMMIO_p = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  toggle_5923_valid_reg = _RAND_100[0:0];
  _RAND_101 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_0_p = _RAND_101[63:0];
  _RAND_102 = {2{`RANDOM}};
  toggle_5924_valid_reg = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_1_p = _RAND_103[63:0];
  _RAND_104 = {2{`RANDOM}};
  toggle_5988_valid_reg = _RAND_104[63:0];
  _RAND_105 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_2_p = _RAND_105[63:0];
  _RAND_106 = {2{`RANDOM}};
  toggle_6052_valid_reg = _RAND_106[63:0];
  _RAND_107 = {2{`RANDOM}};
  wbu_io_in_bits_r_commits_3_p = _RAND_107[63:0];
  _RAND_108 = {2{`RANDOM}};
  toggle_6116_valid_reg = _RAND_108[63:0];
  _RAND_109 = {1{`RANDOM}};
  wbu_io_in_bits_r_isExit_p = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  toggle_6180_valid_reg = _RAND_110[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(valid_t); // @[src/main/scala/utils/Pipeline.scala 24:24]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[5]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[6]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[7]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[8]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[9]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[10]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[11]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[12]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[13]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[14]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[15]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[16]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[17]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[18]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[19]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[20]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[21]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[22]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[23]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[24]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[25]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[26]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[27]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[28]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[29]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[30]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[31]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[32]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[33]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[34]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[35]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[36]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[37]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[38]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[39]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[40]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[41]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[42]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[43]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[44]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[45]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[46]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[47]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[48]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[49]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[50]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[51]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[52]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[53]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[54]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[55]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[56]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[57]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[58]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[59]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[60]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[61]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[62]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_instr_t[63]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[5]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[6]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[7]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[8]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[9]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[10]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[11]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[12]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[13]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[14]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[15]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[16]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[17]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[18]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[19]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[20]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[21]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[22]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[23]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[24]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[25]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[26]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[27]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[28]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[29]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[30]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[31]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[32]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[33]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[34]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[35]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[36]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[37]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pc_t[38]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[5]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[6]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[7]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[8]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[9]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[10]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[11]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[12]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[13]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[14]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[15]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[16]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[17]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[18]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[19]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[20]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[21]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[22]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[23]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[24]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[25]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[26]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[27]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[28]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[29]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[30]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[31]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[32]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[33]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[34]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[35]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[36]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[37]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_pnpc_t[38]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_exceptionVec_1_t); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_exceptionVec_2_t); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_exceptionVec_12_t); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_intrVec_1_t); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_intrVec_3_t); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_intrVec_5_t); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_intrVec_7_t); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_intrVec_9_t); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_intrVec_11_t); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_brIdx_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_brIdx_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_brIdx_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_brIdx_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_cf_crossBoundaryFault_t); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_ctrl_fuType_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_ctrl_fuType_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_ctrl_fuType_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_ctrl_fuOpType_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_ctrl_fuOpType_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_ctrl_fuOpType_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_ctrl_fuOpType_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_ctrl_fuOpType_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_ctrl_fuOpType_t[5]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_ctrl_fuOpType_t[6]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_ctrl_rfWen_t); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_ctrl_rfDest_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_ctrl_rfDest_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_ctrl_rfDest_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_ctrl_rfDest_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_ctrl_rfDest_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_ctrl_isNutCoreTrap_t); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[5]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[6]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[7]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[8]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[9]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[10]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[11]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[12]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[13]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[14]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[15]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[16]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[17]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[18]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[19]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[20]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[21]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[22]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[23]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[24]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[25]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[26]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[27]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[28]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[29]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[30]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[31]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[32]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[33]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[34]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[35]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[36]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[37]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[38]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[39]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[40]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[41]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[42]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[43]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[44]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[45]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[46]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[47]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[48]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[49]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[50]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[51]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[52]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[53]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[54]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[55]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[56]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[57]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[58]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[59]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[60]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[61]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[62]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src1_t[63]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[5]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[6]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[7]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[8]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[9]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[10]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[11]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[12]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[13]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[14]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[15]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[16]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[17]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[18]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[19]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[20]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[21]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[22]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[23]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[24]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[25]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[26]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[27]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[28]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[29]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[30]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[31]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[32]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[33]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[34]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[35]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[36]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[37]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[38]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[39]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[40]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[41]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[42]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[43]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[44]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[45]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[46]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[47]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[48]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[49]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[50]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[51]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[52]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[53]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[54]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[55]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[56]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[57]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[58]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[59]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[60]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[61]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[62]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_src2_t[63]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[5]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[6]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[7]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[8]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[9]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[10]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[11]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[12]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[13]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[14]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[15]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[16]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[17]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[18]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[19]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[20]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[21]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[22]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[23]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[24]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[25]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[26]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[27]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[28]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[29]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[30]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[31]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[32]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[33]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[34]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[35]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[36]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[37]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[38]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[39]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[40]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[41]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[42]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[43]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[44]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[45]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[46]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[47]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[48]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[49]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[50]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[51]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[52]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[53]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[54]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[55]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[56]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[57]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[58]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[59]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[60]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[61]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[62]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(exu_io_in_bits_r_data_imm_t[63]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(valid_1_t); // @[src/main/scala/utils/Pipeline.scala 24:24]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[5]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[6]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[7]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[8]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[9]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[10]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[11]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[12]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[13]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[14]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[15]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[16]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[17]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[18]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[19]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[20]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[21]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[22]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[23]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[24]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[25]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[26]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[27]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[28]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[29]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[30]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[31]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[32]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[33]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[34]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[35]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[36]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[37]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[38]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[39]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[40]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[41]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[42]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[43]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[44]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[45]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[46]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[47]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[48]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[49]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[50]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[51]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[52]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[53]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[54]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[55]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[56]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[57]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[58]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[59]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[60]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[61]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[62]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_instr_t[63]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[5]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[6]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[7]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[8]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[9]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[10]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[11]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[12]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[13]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[14]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[15]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[16]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[17]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[18]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[19]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[20]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[21]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[22]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[23]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[24]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[25]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[26]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[27]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[28]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[29]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[30]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[31]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[32]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[33]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[34]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[35]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[36]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[37]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_pc_t[38]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[5]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[6]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[7]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[8]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[9]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[10]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[11]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[12]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[13]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[14]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[15]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[16]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[17]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[18]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[19]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[20]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[21]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[22]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[23]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[24]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[25]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[26]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[27]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[28]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[29]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[30]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[31]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[32]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[33]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[34]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[35]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[36]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[37]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_target_t[38]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_cf_redirect_valid_t); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_ctrl_fuType_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_ctrl_fuType_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_ctrl_fuType_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_ctrl_rfWen_t); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_ctrl_rfDest_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_ctrl_rfDest_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_ctrl_rfDest_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_ctrl_rfDest_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_decode_ctrl_rfDest_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_isMMIO_t); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[5]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[6]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[7]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[8]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[9]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[10]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[11]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[12]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[13]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[14]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[15]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[16]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[17]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[18]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[19]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[20]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[21]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[22]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[23]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[24]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[25]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[26]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[27]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[28]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[29]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[30]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[31]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[32]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[33]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[34]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[35]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[36]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[37]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[38]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[39]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[40]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[41]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[42]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[43]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[44]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[45]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[46]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[47]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[48]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[49]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[50]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[51]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[52]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[53]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[54]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[55]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[56]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[57]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[58]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[59]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[60]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[61]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[62]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_0_t[63]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[5]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[6]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[7]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[8]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[9]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[10]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[11]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[12]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[13]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[14]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[15]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[16]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[17]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[18]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[19]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[20]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[21]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[22]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[23]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[24]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[25]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[26]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[27]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[28]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[29]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[30]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[31]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[32]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[33]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[34]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[35]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[36]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[37]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[38]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[39]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[40]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[41]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[42]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[43]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[44]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[45]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[46]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[47]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[48]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[49]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[50]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[51]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[52]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[53]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[54]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[55]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[56]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[57]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[58]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[59]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[60]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[61]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[62]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_1_t[63]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[5]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[6]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[7]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[8]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[9]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[10]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[11]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[12]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[13]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[14]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[15]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[16]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[17]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[18]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[19]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[20]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[21]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[22]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[23]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[24]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[25]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[26]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[27]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[28]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[29]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[30]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[31]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[32]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[33]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[34]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[35]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[36]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[37]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[38]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[39]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[40]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[41]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[42]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[43]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[44]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[45]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[46]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[47]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[48]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[49]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[50]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[51]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[52]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[53]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[54]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[55]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[56]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[57]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[58]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[59]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[60]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[61]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[62]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_2_t[63]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[5]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[6]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[7]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[8]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[9]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[10]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[11]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[12]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[13]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[14]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[15]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[16]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[17]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[18]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[19]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[20]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[21]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[22]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[23]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[24]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[25]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[26]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[27]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[28]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[29]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[30]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[31]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[32]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[33]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[34]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[35]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[36]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[37]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[38]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[39]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[40]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[41]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[42]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[43]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[44]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[45]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[46]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[47]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[48]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[49]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[50]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[51]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[52]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[53]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[54]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[55]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[56]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[57]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[58]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[59]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[60]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[61]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[62]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_commits_3_t[63]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(wbu_io_in_bits_r_isExit_t); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
  end
endmodule
module LockingArbiter(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_0_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_in_1_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_1_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_1_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_1_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [7:0]  io_in_1_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_1_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_out_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [7:0]  io_out_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [63:0] io_out_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_chosen // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] lockCount_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  lockIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
  wire  locked = lockCount_value != 3'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 61:34]
  wire  wantsLock = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:62]
  wire  _T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _value_T_1 = lockCount_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  io_chosen_choice = io_in_0_valid ? 1'h0 : 1'h1; // @[src/main/scala/chisel3/util/Arbiter.scala 103:{26,35} 101:41]
  wire  _T_2 = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  wire  _io_in_0_ready_T_1 = locked ? ~lockIdx : 1'h1; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  _io_in_1_ready_T_1 = locked ? lockIdx : _T_2; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [2:0] lockCount_value_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [2:0] lockCount_value_t = lockCount_value ^ lockCount_value_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  toggle_6181_clock;
  wire  toggle_6181_reset;
  wire [2:0] toggle_6181_valid;
  reg [2:0] toggle_6181_valid_reg;
  reg  lockIdx_p; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
  wire  lockIdx_t = lockIdx ^ lockIdx_p; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
  wire  toggle_6184_clock;
  wire  toggle_6184_reset;
  wire  toggle_6184_valid;
  reg  toggle_6184_valid_reg;
  GEN_w3_toggle #(.COVER_INDEX(6181)) toggle_6181 (
    .clock(toggle_6181_clock),
    .reset(toggle_6181_reset),
    .valid(toggle_6181_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(6184)) toggle_6184 (
    .clock(toggle_6184_clock),
    .reset(toggle_6184_reset),
    .valid(toggle_6184_valid)
  );
  assign io_in_0_ready = _io_in_0_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_in_1_ready = _io_in_1_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  assign io_out_bits_addr = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_cmd = io_chosen ? io_in_1_bits_cmd : 4'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wmask = io_chosen ? io_in_1_bits_wmask : 8'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wdata = io_chosen ? io_in_1_bits_wdata : 64'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_chosen = locked ? lockIdx : io_chosen_choice; // @[src/main/scala/chisel3/util/Arbiter.scala 54:13 69:{18,30}]
  assign toggle_6181_clock = clock;
  assign toggle_6181_reset = reset;
  assign toggle_6181_valid = lockCount_value ^ toggle_6181_valid_reg;
  assign toggle_6184_clock = clock;
  assign toggle_6184_reset = reset;
  assign toggle_6184_valid = lockIdx ^ toggle_6184_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      lockCount_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockCount_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockIdx <= io_chosen; // @[src/main/scala/chisel3/util/Arbiter.scala 65:15]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    lockCount_value_p <= lockCount_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    toggle_6181_valid_reg <= lockCount_value;
    lockIdx_p <= lockIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
    toggle_6184_valid_reg <= lockIdx;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lockCount_value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  lockIdx = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  lockCount_value_p = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  toggle_6181_valid_reg = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  lockIdx_p = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  toggle_6184_valid_reg = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(lockCount_value_t[0]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(lockCount_value_t[1]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(lockCount_value_t[2]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(lockIdx_t); // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
    end
  end
endmodule
module SimpleBusCrossbarNto1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_0_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_0_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_0_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_0_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_1_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_1_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_1_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_in_1_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [7:0]  io_in_1_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_in_1_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_1_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_in_1_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_1_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_out_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_out_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_out_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_out_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_out_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_out_resp_bits_rdata // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_reset; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_0_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_1_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_in_1_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_out_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_out_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  reg [1:0] state; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
  wire  _T_1 = ~inputArb_io_out_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:18]
  wire  _T_4 = ~inputArb_io_out_bits_cmd[0] & ~inputArb_io_out_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  reg  inflightSrc; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
  wire  _io_out_req_valid_T = state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 103:47]
  wire  _T_15 = inputArb_io_out_ready & inputArb_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_21 = inputArb_io_out_bits_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire  _T_22 = inputArb_io_out_bits_cmd == 4'h1; // @[src/main/scala/bus/simplebus/SimpleBus.scala 77:29]
  wire [1:0] _GEN_4 = _T_21 | _T_22 ? 2'h2 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 118:{80,88} 92:22]
  wire  _T_25 = io_out_resp_ready & io_out_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_26 = io_out_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:26]
  wire [1:0] _GEN_9 = _T_25 ? 2'h0 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 122:{50,58} 92:22]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [1:0] state_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
  wire [1:0] state_t = state ^ state_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
  wire  toggle_6185_clock;
  wire  toggle_6185_reset;
  wire [1:0] toggle_6185_valid;
  reg [1:0] toggle_6185_valid_reg;
  reg  inflightSrc_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
  wire  inflightSrc_t = inflightSrc ^ inflightSrc_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
  wire  toggle_6187_clock;
  wire  toggle_6187_reset;
  wire  toggle_6187_valid;
  reg  toggle_6187_valid_reg;
  LockingArbiter inputArb ( // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(inputArb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  GEN_w2_toggle #(.COVER_INDEX(6185)) toggle_6185 (
    .clock(toggle_6185_clock),
    .reset(toggle_6185_reset),
    .valid(toggle_6185_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(6187)) toggle_6187 (
    .clock(toggle_6187_clock),
    .reset(toggle_6187_reset),
    .valid(toggle_6187_valid)
  );
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_0_resp_valid = ~inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_1_resp_valid = inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_1_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_out_req_valid = inputArb_io_out_valid & state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 103:37]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_resp_ready = 1'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 110:{13,13}]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_wmask = io_in_1_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_out_ready = io_out_req_ready & _io_out_req_valid_T; // @[src/main/scala/bus/simplebus/Crossbar.scala 104:37]
  assign toggle_6185_clock = clock;
  assign toggle_6185_reset = reset;
  assign toggle_6185_valid = state ^ toggle_6185_valid_reg;
  assign toggle_6187_clock = clock;
  assign toggle_6187_reset = reset;
  assign toggle_6187_valid = inflightSrc ^ toggle_6187_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
      state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_15) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:29]
        if (_T_4) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 117:38]
          state <= 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 117:46]
        end else begin
          state <= _GEN_4;
        end
      end
    end else if (2'h1 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_25 & _T_26) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 121:82]
        state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 121:90]
      end
    end else if (2'h2 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      state <= _GEN_9;
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
      inflightSrc <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_15) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:29]
        inflightSrc <= inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 116:21]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(inputArb_io_out_valid & ~_T_4 & _T_1))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Crossbar.scala:98 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"
            ); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    state_p <= state; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
    toggle_6185_valid_reg <= state;
    inflightSrc_p <= inflightSrc; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
    toggle_6187_valid_reg <= inflightSrc;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  inflightSrc = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_p = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  toggle_6185_valid_reg = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  inflightSrc_p = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  toggle_6187_valid_reg = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~(inputArb_io_out_valid & ~_T_4 & _T_1)); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
    end
    //
    if (enToggle_past) begin
      cover(state_t[0]); // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[1]); // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
    end
    //
    if (enToggle_past) begin
      cover(inflightSrc_t); // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
    end
  end
endmodule
module LockingArbiter_1(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_0_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [2:0]  io_in_0_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_0_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [7:0]  io_in_0_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_0_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_in_1_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_1_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_1_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_1_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_1_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_in_2_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_2_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_2_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_2_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_2_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_out_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [2:0]  io_out_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [7:0]  io_out_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [63:0] io_out_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [1:0]  io_chosen // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  _GEN_1 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  wire  _GEN_2 = 2'h2 == io_chosen ? io_in_2_valid : _GEN_1; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  wire [31:0] _GEN_5 = 2'h1 == io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [31:0] _GEN_6 = 2'h2 == io_chosen ? io_in_2_bits_addr : _GEN_5; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [2:0] _GEN_9 = 2'h1 == io_chosen ? 3'h3 : io_in_0_bits_size; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [2:0] _GEN_10 = 2'h2 == io_chosen ? 3'h3 : _GEN_9; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [3:0] _GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_cmd : io_in_0_bits_cmd; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [3:0] _GEN_14 = 2'h2 == io_chosen ? io_in_2_bits_cmd : _GEN_13; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [7:0] _GEN_17 = 2'h1 == io_chosen ? 8'hff : io_in_0_bits_wmask; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [7:0] _GEN_18 = 2'h2 == io_chosen ? 8'hff : _GEN_17; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [63:0] _GEN_21 = 2'h1 == io_chosen ? io_in_1_bits_wdata : io_in_0_bits_wdata; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  wire [63:0] _GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_wdata : _GEN_21; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  reg [2:0] lockCount_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [1:0] lockIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
  wire  locked = lockCount_value != 3'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 61:34]
  wire  wantsLock = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:62]
  wire  _T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _value_T_1 = lockCount_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [1:0] _GEN_27 = io_in_2_valid ? 2'h2 : 2'h3; // @[src/main/scala/chisel3/util/Arbiter.scala 103:{26,35} 101:41]
  wire [1:0] _GEN_28 = io_in_1_valid ? 2'h1 : _GEN_27; // @[src/main/scala/chisel3/util/Arbiter.scala 103:{26,35}]
  wire [1:0] io_chosen_choice = io_in_0_valid ? 2'h0 : _GEN_28; // @[src/main/scala/chisel3/util/Arbiter.scala 103:{26,35}]
  wire  _T_4 = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  wire  _T_5 = ~(io_in_0_valid | io_in_1_valid); // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  wire  _io_in_0_ready_T_1 = locked ? lockIdx == 2'h0 : 1'h1; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  _io_in_1_ready_T_1 = locked ? lockIdx == 2'h1 : _T_4; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  _io_in_2_ready_T_1 = locked ? lockIdx == 2'h2 : _T_5; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [2:0] lockCount_value_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [2:0] lockCount_value_t = lockCount_value ^ lockCount_value_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  toggle_6188_clock;
  wire  toggle_6188_reset;
  wire [2:0] toggle_6188_valid;
  reg [2:0] toggle_6188_valid_reg;
  reg [1:0] lockIdx_p; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
  wire [1:0] lockIdx_t = lockIdx ^ lockIdx_p; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
  wire  toggle_6191_clock;
  wire  toggle_6191_reset;
  wire [1:0] toggle_6191_valid;
  reg [1:0] toggle_6191_valid_reg;
  GEN_w3_toggle #(.COVER_INDEX(6188)) toggle_6188 (
    .clock(toggle_6188_clock),
    .reset(toggle_6188_reset),
    .valid(toggle_6188_valid)
  );
  GEN_w2_toggle #(.COVER_INDEX(6191)) toggle_6191 (
    .clock(toggle_6191_clock),
    .reset(toggle_6191_reset),
    .valid(toggle_6191_valid)
  );
  assign io_in_0_ready = _io_in_0_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_in_1_ready = _io_in_1_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_in_2_ready = _io_in_2_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_out_valid = 2'h3 == io_chosen ? 1'h0 : _GEN_2; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  assign io_out_bits_addr = 2'h3 == io_chosen ? 32'h0 : _GEN_6; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_size = 2'h3 == io_chosen ? 3'h0 : _GEN_10; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_cmd = 2'h3 == io_chosen ? 4'h0 : _GEN_14; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wmask = 2'h3 == io_chosen ? 8'h0 : _GEN_18; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wdata = 2'h3 == io_chosen ? 64'h0 : _GEN_22; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_chosen = locked ? lockIdx : io_chosen_choice; // @[src/main/scala/chisel3/util/Arbiter.scala 54:13 69:{18,30}]
  assign toggle_6188_clock = clock;
  assign toggle_6188_reset = reset;
  assign toggle_6188_valid = lockCount_value ^ toggle_6188_valid_reg;
  assign toggle_6191_clock = clock;
  assign toggle_6191_reset = reset;
  assign toggle_6191_valid = lockIdx ^ toggle_6191_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      lockCount_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockCount_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockIdx <= io_chosen; // @[src/main/scala/chisel3/util/Arbiter.scala 65:15]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    lockCount_value_p <= lockCount_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    toggle_6188_valid_reg <= lockCount_value;
    lockIdx_p <= lockIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
    toggle_6191_valid_reg <= lockIdx;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lockCount_value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  lockIdx = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  lockCount_value_p = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  toggle_6188_valid_reg = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  lockIdx_p = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  toggle_6191_valid_reg = _RAND_5[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(lockCount_value_t[0]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(lockCount_value_t[1]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(lockCount_value_t[2]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(lockIdx_t[0]); // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
    end
    //
    if (enToggle_past) begin
      cover(lockIdx_t[1]); // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
    end
  end
endmodule
module SimpleBusCrossbarNto1_1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_0_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_0_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [2:0]  io_in_0_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_in_0_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [7:0]  io_in_0_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_in_0_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_0_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_0_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_1_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_1_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_1_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_in_1_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_in_1_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_1_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_1_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_2_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_2_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_2_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_in_2_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_in_2_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_2_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_2_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_out_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_out_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [2:0]  io_out_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_out_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_out_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_out_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_out_resp_bits_rdata // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_reset; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_0_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [2:0] inputArb_io_in_0_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_0_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_in_0_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_0_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_1_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_2_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_2_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_2_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_2_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_2_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_out_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_out_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [2:0] inputArb_io_out_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [1:0] inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  reg [1:0] state; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
  wire  _T_1 = ~inputArb_io_out_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:18]
  wire  _T_4 = ~inputArb_io_out_bits_cmd[0] & ~inputArb_io_out_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  reg [1:0] inflightSrc; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
  wire  _io_out_req_valid_T = state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 103:47]
  wire  _T_15 = inputArb_io_out_ready & inputArb_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_21 = inputArb_io_out_bits_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire  _T_22 = inputArb_io_out_bits_cmd == 4'h1; // @[src/main/scala/bus/simplebus/SimpleBus.scala 77:29]
  wire [1:0] _GEN_8 = _T_21 | _T_22 ? 2'h2 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 118:{80,88} 92:22]
  wire  _T_25 = io_out_resp_ready & io_out_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_26 = io_out_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:26]
  wire [1:0] _GEN_13 = _T_25 ? 2'h0 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 122:{50,58} 92:22]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [1:0] state_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
  wire [1:0] state_t = state ^ state_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
  wire  toggle_6193_clock;
  wire  toggle_6193_reset;
  wire [1:0] toggle_6193_valid;
  reg [1:0] toggle_6193_valid_reg;
  reg [1:0] inflightSrc_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
  wire [1:0] inflightSrc_t = inflightSrc ^ inflightSrc_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
  wire  toggle_6195_clock;
  wire  toggle_6195_reset;
  wire [1:0] toggle_6195_valid;
  reg [1:0] toggle_6195_valid_reg;
  LockingArbiter_1 inputArb ( // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_0_bits_size(inputArb_io_in_0_bits_size),
    .io_in_0_bits_cmd(inputArb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(inputArb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(inputArb_io_in_0_bits_wdata),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_in_2_ready(inputArb_io_in_2_ready),
    .io_in_2_valid(inputArb_io_in_2_valid),
    .io_in_2_bits_addr(inputArb_io_in_2_bits_addr),
    .io_in_2_bits_cmd(inputArb_io_in_2_bits_cmd),
    .io_in_2_bits_wdata(inputArb_io_in_2_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_size(inputArb_io_out_bits_size),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  GEN_w2_toggle #(.COVER_INDEX(6193)) toggle_6193 (
    .clock(toggle_6193_clock),
    .reset(toggle_6193_reset),
    .valid(toggle_6193_valid)
  );
  GEN_w2_toggle #(.COVER_INDEX(6195)) toggle_6195 (
    .clock(toggle_6195_clock),
    .reset(toggle_6195_reset),
    .valid(toggle_6195_valid)
  );
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_0_resp_valid = 2'h0 == inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_1_resp_valid = 2'h1 == inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_2_req_ready = inputArb_io_in_2_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_2_resp_valid = 2'h2 == inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_2_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_out_req_valid = inputArb_io_out_valid & state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 103:37]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_size = inputArb_io_out_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_resp_ready = 1'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 110:{13,13}]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_size = io_in_0_req_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_cmd = io_in_0_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_wmask = io_in_0_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_2_valid = io_in_2_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_2_bits_addr = io_in_2_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_2_bits_cmd = io_in_2_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_2_bits_wdata = io_in_2_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_out_ready = io_out_req_ready & _io_out_req_valid_T; // @[src/main/scala/bus/simplebus/Crossbar.scala 104:37]
  assign toggle_6193_clock = clock;
  assign toggle_6193_reset = reset;
  assign toggle_6193_valid = state ^ toggle_6193_valid_reg;
  assign toggle_6195_clock = clock;
  assign toggle_6195_reset = reset;
  assign toggle_6195_valid = inflightSrc ^ toggle_6195_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
      state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_15) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:29]
        if (_T_4) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 117:38]
          state <= 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 117:46]
        end else begin
          state <= _GEN_8;
        end
      end
    end else if (2'h1 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_25 & _T_26) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 121:82]
        state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 121:90]
      end
    end else if (2'h2 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      state <= _GEN_13;
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
      inflightSrc <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_15) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:29]
        inflightSrc <= inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 116:21]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(inputArb_io_out_valid & ~_T_4 & _T_1))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Crossbar.scala:98 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"
            ); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    state_p <= state; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
    toggle_6193_valid_reg <= state;
    inflightSrc_p <= inflightSrc; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
    toggle_6195_valid_reg <= inflightSrc;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  inflightSrc = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  state_p = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  toggle_6193_valid_reg = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  inflightSrc_p = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  toggle_6195_valid_reg = _RAND_5[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~(inputArb_io_out_valid & ~_T_4 & _T_1)); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
    end
    //
    if (enToggle_past) begin
      cover(state_t[0]); // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[1]); // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
    end
    //
    if (enToggle_past) begin
      cover(inflightSrc_t[0]); // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
    end
    //
    if (enToggle_past) begin
      cover(inflightSrc_t[1]); // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
    end
  end
endmodule
module EmbeddedTLBExec(
  input          clock,
  input          reset,
  output         io_in_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_in_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [38:0]  io_in_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [86:0]  io_in_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_out_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_out_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [31:0]  io_out_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [86:0]  io_out_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_0, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_1, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_2, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_3, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_mdWrite_wen, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [3:0]   io_mdWrite_waymask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [144:0] io_mdWrite_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_mdReady, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_mem_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_mem_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [31:0]  io_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [3:0]   io_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [63:0]  io_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_mem_resp_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_mem_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [63:0]  io_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_flush, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [63:0]  io_satp, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [1:0]   io_pf_priviledgeMode, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_loadPF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_storePF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_laf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_saf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_ipf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_iaf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_isFinish // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] vpn_vpn0 = io_in_bits_addr[20:12]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:54]
  wire [8:0] vpn_vpn1 = io_in_bits_addr[29:21]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:54]
  wire [8:0] vpn_vpn2 = io_in_bits_addr[38:30]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:54]
  wire [43:0] satp_ppn = io_satp[43:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 244:30]
  wire [15:0] satp_asid = io_satp[59:44]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 244:30]
  wire [17:0] hitVec_hi = {vpn_vpn2,vpn_vpn1}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:201]
  wire [26:0] _hitVec_T_34 = {vpn_vpn2,vpn_vpn1,vpn_vpn0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:201]
  wire [26:0] _hitVec_T_35 = {9'h1ff,io_md_0[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_36 = _hitVec_T_35 & io_md_0[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_38 = _hitVec_T_35 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_39 = _hitVec_T_36 == _hitVec_T_38; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_40 = io_md_0[76] & io_md_0[117:102] == satp_asid & _hitVec_T_39; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [26:0] _hitVec_T_76 = {9'h1ff,io_md_1[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_77 = _hitVec_T_76 & io_md_1[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_79 = _hitVec_T_76 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_80 = _hitVec_T_77 == _hitVec_T_79; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_81 = io_md_1[76] & io_md_1[117:102] == satp_asid & _hitVec_T_80; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [26:0] _hitVec_T_117 = {9'h1ff,io_md_2[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_118 = _hitVec_T_117 & io_md_2[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_120 = _hitVec_T_117 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_121 = _hitVec_T_118 == _hitVec_T_120; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_122 = io_md_2[76] & io_md_2[117:102] == satp_asid & _hitVec_T_121; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [26:0] _hitVec_T_158 = {9'h1ff,io_md_3[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_159 = _hitVec_T_158 & io_md_3[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_161 = _hitVec_T_158 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_162 = _hitVec_T_159 == _hitVec_T_161; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_163 = io_md_3[76] & io_md_3[117:102] == satp_asid & _hitVec_T_162; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [3:0] hitVec = {_hitVec_T_163,_hitVec_T_122,_hitVec_T_81,_hitVec_T_40}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:211]
  wire  _hit_T = |hitVec; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 249:35]
  wire  hit = io_in_valid & |hitVec; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 249:25]
  wire  miss = io_in_valid & ~_hit_T; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 250:26]
  reg [63:0] victimWaymask_lfsr; // @[src/main/scala/utils/LFSR64.scala 25:23]
  wire  victimWaymask_xor = victimWaymask_lfsr[0] ^ victimWaymask_lfsr[1] ^ victimWaymask_lfsr[3] ^ victimWaymask_lfsr[4
    ]; // @[src/main/scala/utils/LFSR64.scala 26:43]
  wire [63:0] _victimWaymask_lfsr_T_2 = {victimWaymask_xor,victimWaymask_lfsr[63:1]}; // @[src/main/scala/utils/LFSR64.scala 28:41]
  wire [3:0] victimWaymask = 4'h1 << victimWaymask_lfsr[1:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 252:42]
  wire [3:0] waymask = hit ? hitVec : victimWaymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:20]
  wire [144:0] _hitMeta_T_4 = waymask[0] ? io_md_0 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_5 = waymask[1] ? io_md_1 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_6 = waymask[2] ? io_md_2 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_7 = waymask[3] ? io_md_3 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_8 = _hitMeta_T_4 | _hitMeta_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_9 = _hitMeta_T_8 | _hitMeta_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_10 = _hitMeta_T_9 | _hitMeta_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] hitMeta_flag = _hitMeta_T_10[83:76]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 262:70]
  wire [17:0] hitMeta_mask = _hitMeta_T_10[101:84]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 262:70]
  wire [43:0] hitData_ppn = _hitMeta_T_10[75:32]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 263:70]
  wire  hitFlag_x = hitMeta_flag[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_u = hitMeta_flag[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_a = hitMeta_flag[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  _hitCheck_T = io_pf_priviledgeMode == 2'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:62]
  wire  _hitCheck_T_5 = io_pf_priviledgeMode == 2'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:110]
  wire  hitCheck = hit & ~(io_pf_priviledgeMode == 2'h0 & ~hitFlag_u) & ~(io_pf_priviledgeMode == 2'h1 & hitFlag_u); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:87]
  wire  hitADCheck = ~hitFlag_a; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 274:20]
  wire  hitExec = hitCheck & ~hitADCheck & hitFlag_x; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:41]
  wire  hitinstrPF = ~hitExec & hit; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 290:52]
  reg [2:0] state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
  reg [1:0] level; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
  reg [63:0] memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
  reg [17:0] missMaskStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
  wire  memRdata_flag_v = io_mem_resp_bits_rdata[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_r = io_mem_resp_bits_rdata[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_w = io_mem_resp_bits_rdata[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_x = io_mem_resp_bits_rdata[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_u = io_mem_resp_bits_rdata[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_g = io_mem_resp_bits_rdata[5]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_a = io_mem_resp_bits_rdata[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_d = io_mem_resp_bits_rdata[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire [43:0] memRdata_ppn = io_mem_resp_bits_rdata[53:10]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire [9:0] memRdata_reserved = io_mem_resp_bits_rdata[63:54]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  reg [55:0] raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
  wire  _raddrCancel_T_3 = |(raddr >= 56'h80000000 & raddr < 56'h100000000); // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  raddrCancel = ~_raddrCancel_T_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 308:21]
  wire  _alreadyOutFire_T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  alreadyOutFire; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
  wire  _GEN_2 = _alreadyOutFire_T | alreadyOutFire; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:{33,33,33}]
  reg  needFlush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 312:26]
  wire  isFlush = needFlush | io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 314:27]
  wire  _GEN_3 = io_flush & state != 3'h0 | needFlush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 312:26 315:{40,52}]
  wire  _GEN_4 = _alreadyOutFire_T & needFlush ? 1'h0 : _GEN_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 316:{37,49}]
  reg  missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24]
  reg  missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
  wire  _T_5 = ~io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 324:13]
  wire [55:0] _raddr_T_1 = {satp_ppn,vpn_vpn2,3'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 89:8]
  wire  _T_10 = io_mem_req_ready & io_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _GEN_15 = raddrCancel ? 3'h4 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 343:32 344:29]
  wire  _GEN_16 = raddrCancel | missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 343:32 345:19 319:26]
  wire [2:0] _GEN_17 = _T_10 ? 3'h2 : _GEN_15; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 341:38 342:15]
  wire  _GEN_18 = _T_10 ? missPTEAF : _GEN_16; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26 341:38]
  wire  _GEN_20 = isFlush ? 1'h0 : _GEN_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 338:22 340:19]
  wire [7:0] _missflag_T = {memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,memRdata_flag_u,memRdata_flag_x,
    memRdata_flag_w,memRdata_flag_r,memRdata_flag_v}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_v = _missflag_T[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_r = _missflag_T[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_w = _missflag_T[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_x = _missflag_T[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_u = _missflag_T[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_g = _missflag_T[5]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_a = _missflag_T[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_d = _missflag_T[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  _T_12 = io_mem_resp_ready & io_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_15 = level == 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:58]
  wire  _T_16 = level == 2'h2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:73]
  wire  _T_21 = ~missflag_r & missflag_w; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:44]
  wire [8:0] _raddr_T_3 = _T_15 ? vpn_vpn1 : vpn_vpn0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 369:50]
  wire [55:0] _raddr_T_5 = {memRdata_ppn,_raddr_T_3,3'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 89:8]
  wire  is_reserved = memRdata_reserved != 10'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 370:49]
  wire [2:0] _GEN_22 = is_reserved ? 3'h4 : 3'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 368:19 371:32 372:21]
  wire  _GEN_23 = is_reserved | missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24 371:32 374:25]
  wire [2:0] _GEN_24 = ~missflag_v | ~missflag_r & missflag_w ? 3'h4 : _GEN_22; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:60 357:43]
  wire  _GEN_25 = ~missflag_v | ~missflag_r & missflag_w | _GEN_23; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:60 358:45]
  wire [55:0] _GEN_26 = ~missflag_v | ~missflag_r & missflag_w ? raddr : _raddr_T_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18 356:60 369:19]
  wire [17:0] pg_mask = _T_16 ? 18'h1ff : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 384:28]
  wire [43:0] _GEN_121 = {{26'd0}, pg_mask}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:54]
  wire [43:0] _misaligned_T_1 = memRdata_ppn & _GEN_121; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:54]
  wire  misaligned = level[1] & |_misaligned_T_1 | is_reserved; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:76]
  wire  permCheck = missflag_v & ~(_hitCheck_T & ~missflag_u) & ~(_hitCheck_T_5 & missflag_u); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 386:87]
  wire  permAD = ~missflag_a; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 388:24]
  wire  permExec = permCheck & ~_T_21 & ~permAD & ~misaligned & missflag_x; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 389:75]
  wire [7:0] _missRefillFlag_T_2 = {missflag_d,missflag_a,missflag_g,missflag_u,missflag_x,missflag_w,missflag_r,
    missflag_v}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 393:79]
  wire [7:0] _missRefillFlag_T_3 = 8'h40 | _missRefillFlag_T_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 393:68]
  wire [63:0] _memRespStore_T = io_mem_resp_bits_rdata | 64'h40; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 394:50]
  wire  _GEN_27 = ~permExec | missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24 396:{30,40}]
  wire  _GEN_29 = ~permExec ? 1'h0 : 1'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 396:30 304:32 399:30]
  wire [17:0] _missMask_T_2 = _T_16 ? 18'h3fe00 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 412:59]
  wire [17:0] _missMask_T_3 = _T_15 ? 18'h0 : _missMask_T_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 412:26]
  wire [7:0] _GEN_30 = level != 2'h0 ? _missRefillFlag_T_3 : 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 393:26 305:32]
  wire [63:0] _GEN_31 = level != 2'h0 ? _memRespStore_T : memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 394:24 301:25]
  wire  _GEN_32 = level != 2'h0 ? _GEN_27 : missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24 383:36]
  wire [2:0] _GEN_33 = level != 2'h0 ? 3'h4 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 383:36]
  wire  _GEN_34 = level != 2'h0 & _GEN_29; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 383:36]
  wire [17:0] _GEN_35 = level != 2'h0 ? _missMask_T_3 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 412:20 302:26]
  wire [17:0] _GEN_43 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 18'h3ffff : _GEN_35; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26 355:82]
  wire [17:0] _GEN_51 = isFlush ? 18'h3ffff : _GEN_43; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 352:24 302:26]
  wire [17:0] _GEN_60 = _T_12 ? _GEN_51 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26 351:33]
  wire [17:0] _GEN_87 = 3'h2 == state ? _GEN_60 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 302:26]
  wire [17:0] _GEN_100 = 3'h1 == state ? 18'h3ffff : _GEN_87; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 302:26]
  wire [17:0] missMask = 3'h0 == state ? 18'h3ffff : _GEN_100; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 302:26]
  wire [17:0] _GEN_36 = level != 2'h0 ? missMask : missMaskStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 413:25 303:26]
  wire [2:0] _GEN_37 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_24 : _GEN_33; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:82]
  wire  _GEN_38 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_25 : _GEN_32; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:82]
  wire [55:0] _GEN_39 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_26 : raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18 355:82]
  wire [7:0] _GEN_40 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 8'h0 : _GEN_30; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32 355:82]
  wire [63:0] _GEN_41 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? memRespStore : _GEN_31; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25 355:82]
  wire  _GEN_42 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 1'h0 : _GEN_34; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 355:82]
  wire [17:0] _GEN_44 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? missMaskStore : _GEN_36; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26 355:82]
  wire [2:0] _GEN_45 = isFlush ? 3'h0 : _GEN_37; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 352:24 353:17]
  wire  _GEN_46 = isFlush ? missIPF : _GEN_38; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24 352:24]
  wire [55:0] _GEN_47 = isFlush ? raddr : _GEN_39; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18 352:24]
  wire [7:0] _GEN_48 = isFlush ? 8'h0 : _GEN_40; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 352:24 305:32]
  wire [63:0] _GEN_49 = isFlush ? memRespStore : _GEN_41; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 352:24 301:25]
  wire  _GEN_50 = isFlush ? 1'h0 : _GEN_42; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 352:24 304:32]
  wire [17:0] _GEN_52 = isFlush ? missMaskStore : _GEN_44; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 352:24 303:26]
  wire [1:0] _level_T_1 = level - 2'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 415:24]
  wire [2:0] _GEN_53 = _T_12 ? _GEN_45 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 351:33]
  wire  _GEN_54 = _T_12 ? _GEN_20 : _GEN_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
  wire  _GEN_55 = _T_12 ? _GEN_46 : missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24 351:33]
  wire  _GEN_59 = _T_12 & _GEN_50; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 351:33]
  wire [1:0] _GEN_62 = _T_12 ? _level_T_1 : level; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33 415:15 299:22]
  wire [2:0] _GEN_63 = _T_10 ? 3'h4 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 423:{38,46}]
  wire [2:0] _GEN_64 = isFlush ? 3'h0 : _GEN_63; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 420:22 421:15]
  wire [2:0] _GEN_65 = io_isFinish | io_flush | alreadyOutFire ? 3'h0 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 427:13 298:22]
  wire  _GEN_66 = io_isFinish | io_flush | alreadyOutFire ? 1'h0 : missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 428:15 318:24]
  wire  _GEN_67 = io_isFinish | io_flush | alreadyOutFire ? 1'h0 : missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 429:17 319:26]
  wire  _GEN_68 = io_isFinish | io_flush | alreadyOutFire ? 1'h0 : _GEN_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 430:22]
  wire [2:0] _GEN_69 = 3'h5 == state ? 3'h0 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 434:13 298:22]
  wire  _GEN_70 = 3'h5 == state ? 1'h0 : missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 435:17 319:26]
  wire [2:0] _GEN_71 = 3'h4 == state ? _GEN_65 : _GEN_69; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_72 = 3'h4 == state ? _GEN_66 : missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 318:24]
  wire  _GEN_73 = 3'h4 == state ? _GEN_67 : _GEN_70; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_74 = 3'h4 == state ? _GEN_68 : _GEN_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire [2:0] _GEN_75 = 3'h3 == state ? _GEN_64 : _GEN_71; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_76 = 3'h3 == state ? _GEN_20 : _GEN_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_77 = 3'h3 == state ? missIPF : _GEN_72; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 318:24]
  wire  _GEN_78 = 3'h3 == state ? missPTEAF : _GEN_73; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 319:26]
  wire  _GEN_79 = 3'h3 == state ? _GEN_2 : _GEN_74; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_99 = 3'h1 == state ? 1'h0 : 3'h2 == state & _GEN_59; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 304:32]
  wire  missMetaRefill = 3'h0 == state ? 1'h0 : _GEN_99; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 304:32]
  wire  cmd = state == 3'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:23]
  wire  _io_mem_req_valid_T_3 = ~isFlush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 442:76]
  wire  _T_34 = missMetaRefill & _io_mem_req_valid_T_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:50]
  wire  _T_35 = state == 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:82]
  reg  REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
  reg [3:0] REG_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:60]
  reg [26:0] REG_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
  reg [15:0] REG_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
  reg [17:0] REG_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
  reg [7:0] REG_6; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
  reg [43:0] REG_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
  reg [55:0] REG_8; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
  wire [168:0] _io_mdWrite_wdata_T = {REG_3,REG_4,REG_5,REG_6,REG_7,REG_8}; // @[src/main/scala/nutcore/mem/TLB.scala 220:22]
  wire [55:0] mdWriteAddr = {memRdata_ppn,12'h0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 451:24]
  wire  _mdMayHasAF_T_2 = mdWriteAddr >= 56'h40000000 & mdWriteAddr < 56'h40001000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_5 = mdWriteAddr >= 56'h80000000 & mdWriteAddr < 56'h100000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [1:0] _mdMayHasAF_T_6 = {_mdMayHasAF_T_5,_mdMayHasAF_T_2}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _mdMayHasAF_T_7 = |_mdMayHasAF_T_6; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  _mdMayHasAF_T_11 = mdWriteAddr >= 56'h38000000 & mdWriteAddr < 56'h38010000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_14 = mdWriteAddr >= 56'h3c000000 & mdWriteAddr < 56'h40000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_17 = mdWriteAddr >= 56'h40600000 & mdWriteAddr < 56'h40600010; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_20 = mdWriteAddr >= 56'h50000000 & mdWriteAddr < 56'h50400000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_23 = mdWriteAddr >= 56'h40001000 & mdWriteAddr < 56'h40001008; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_29 = mdWriteAddr >= 56'h40002000 & mdWriteAddr < 56'h40003000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [7:0] _mdMayHasAF_T_33 = {_mdMayHasAF_T_5,_mdMayHasAF_T_29,_mdMayHasAF_T_2,_mdMayHasAF_T_23,_mdMayHasAF_T_20,
    _mdMayHasAF_T_17,_mdMayHasAF_T_14,_mdMayHasAF_T_11}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _mdMayHasAF_T_34 = |_mdMayHasAF_T_33; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  mdMayHasAF = ~_mdMayHasAF_T_7 | ~_mdMayHasAF_T_34 | ~_mdMayHasAF_T_34; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 452:84]
  reg  blockRefill; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
  wire [55:0] vaddr_ext = {24'h0,io_in_bits_addr[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [55:0] _paddr_T = {hitData_ppn,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:24]
  wire [55:0] _paddr_T_2 = {26'h3ffffff,hitMeta_mask,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:49]
  wire [55:0] _paddr_T_3 = _paddr_T & _paddr_T_2; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [55:0] _paddr_T_4 = ~_paddr_T_2; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [55:0] _paddr_T_5 = vaddr_ext & _paddr_T_4; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [55:0] _paddr_T_6 = _paddr_T_3 | _paddr_T_5; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [55:0] _paddr_T_18 = {memRespStore[53:10],12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:24]
  wire [55:0] _paddr_T_20 = {26'h3ffffff,missMaskStore,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:49]
  wire [55:0] _paddr_T_21 = _paddr_T_18 & _paddr_T_20; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [55:0] _paddr_T_22 = ~_paddr_T_20; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [55:0] _paddr_T_23 = vaddr_ext & _paddr_T_22; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [55:0] _paddr_T_24 = _paddr_T_21 | _paddr_T_23; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [55:0] paddr = hit ? _paddr_T_6 : _paddr_T_24; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 461:15]
  wire  out_req_valid = io_in_valid & (hit | state == 3'h4); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 484:35]
  wire  _instrAF_T_2 = paddr >= 56'h40000000 & paddr < 56'h40001000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _instrAF_T_5 = paddr >= 56'h80000000 & paddr < 56'h100000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [1:0] _instrAF_T_6 = {_instrAF_T_5,_instrAF_T_2}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _instrAF_T_7 = |_instrAF_T_6; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  _hasException_T = io_pf_loadPF | io_pf_storePF; // @[src/main/scala/nutcore/Bundle.scala 134:23]
  wire  _hasException_T_1 = io_pf_laf | io_pf_saf; // @[src/main/scala/nutcore/Bundle.scala 135:24]
  wire  hasException = _hasException_T | _hasException_T_1; // @[src/main/scala/nutcore/Bundle.scala 136:35]
  wire  _io_out_valid_T_5 = ~hasException; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 496:78]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [63:0] victimWaymask_lfsr_p; // @[src/main/scala/utils/LFSR64.scala 25:23]
  wire [63:0] victimWaymask_lfsr_t = victimWaymask_lfsr ^ victimWaymask_lfsr_p; // @[src/main/scala/utils/LFSR64.scala 25:23]
  wire  toggle_6197_clock;
  wire  toggle_6197_reset;
  wire [63:0] toggle_6197_valid;
  reg [63:0] toggle_6197_valid_reg;
  reg [2:0] state_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
  wire [2:0] state_t = state ^ state_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
  wire  toggle_6261_clock;
  wire  toggle_6261_reset;
  wire [2:0] toggle_6261_valid;
  reg [2:0] toggle_6261_valid_reg;
  reg [1:0] level_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
  wire [1:0] level_t = level ^ level_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
  wire  toggle_6264_clock;
  wire  toggle_6264_reset;
  wire [1:0] toggle_6264_valid;
  reg [1:0] toggle_6264_valid_reg;
  reg [63:0] memRespStore_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
  wire [63:0] memRespStore_t = memRespStore ^ memRespStore_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
  wire  toggle_6266_clock;
  wire  toggle_6266_reset;
  wire [63:0] toggle_6266_valid;
  reg [63:0] toggle_6266_valid_reg;
  reg [17:0] missMaskStore_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
  wire [17:0] missMaskStore_t = missMaskStore ^ missMaskStore_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
  wire  toggle_6330_clock;
  wire  toggle_6330_reset;
  wire [17:0] toggle_6330_valid;
  reg [17:0] toggle_6330_valid_reg;
  reg [55:0] raddr_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
  wire [55:0] raddr_t = raddr ^ raddr_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
  wire  toggle_6348_clock;
  wire  toggle_6348_reset;
  wire [55:0] toggle_6348_valid;
  reg [55:0] toggle_6348_valid_reg;
  reg  alreadyOutFire_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
  wire  alreadyOutFire_t = alreadyOutFire ^ alreadyOutFire_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
  wire  toggle_6404_clock;
  wire  toggle_6404_reset;
  wire  toggle_6404_valid;
  reg  toggle_6404_valid_reg;
  reg  needFlush_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 312:26]
  wire  needFlush_t = needFlush ^ needFlush_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 312:26]
  wire  toggle_6405_clock;
  wire  toggle_6405_reset;
  wire  toggle_6405_valid;
  reg  toggle_6405_valid_reg;
  reg  missIPF_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24]
  wire  missIPF_t = missIPF ^ missIPF_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24]
  wire  toggle_6406_clock;
  wire  toggle_6406_reset;
  wire  toggle_6406_valid;
  reg  toggle_6406_valid_reg;
  reg  missPTEAF_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
  wire  missPTEAF_t = missPTEAF ^ missPTEAF_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
  wire  toggle_6407_clock;
  wire  toggle_6407_reset;
  wire  toggle_6407_valid;
  reg  toggle_6407_valid_reg;
  reg  REG_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
  wire  REG_t = REG ^ REG_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
  wire  toggle_6408_clock;
  wire  toggle_6408_reset;
  wire  toggle_6408_valid;
  reg  toggle_6408_valid_reg;
  reg [3:0] REG_2_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:60]
  wire [3:0] REG_2_t = REG_2 ^ REG_2_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:60]
  wire  toggle_6409_clock;
  wire  toggle_6409_reset;
  wire [3:0] toggle_6409_valid;
  reg [3:0] toggle_6409_valid_reg;
  reg [26:0] REG_3_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
  wire [26:0] REG_3_t = REG_3 ^ REG_3_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
  wire  toggle_6413_clock;
  wire  toggle_6413_reset;
  wire [26:0] toggle_6413_valid;
  reg [26:0] toggle_6413_valid_reg;
  reg [15:0] REG_4_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
  wire [15:0] REG_4_t = REG_4 ^ REG_4_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
  wire  toggle_6440_clock;
  wire  toggle_6440_reset;
  wire [15:0] toggle_6440_valid;
  reg [15:0] toggle_6440_valid_reg;
  reg [17:0] REG_5_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
  wire [17:0] REG_5_t = REG_5 ^ REG_5_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
  wire  toggle_6456_clock;
  wire  toggle_6456_reset;
  wire [17:0] toggle_6456_valid;
  reg [17:0] toggle_6456_valid_reg;
  reg [7:0] REG_6_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
  wire [7:0] REG_6_t = REG_6 ^ REG_6_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
  wire  toggle_6474_clock;
  wire  toggle_6474_reset;
  wire [7:0] toggle_6474_valid;
  reg [7:0] toggle_6474_valid_reg;
  reg [43:0] REG_7_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
  wire [43:0] REG_7_t = REG_7 ^ REG_7_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
  wire  toggle_6482_clock;
  wire  toggle_6482_reset;
  wire [43:0] toggle_6482_valid;
  reg [43:0] toggle_6482_valid_reg;
  reg [55:0] REG_8_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
  wire [55:0] REG_8_t = REG_8 ^ REG_8_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
  wire  toggle_6526_clock;
  wire  toggle_6526_reset;
  wire [55:0] toggle_6526_valid;
  reg [55:0] toggle_6526_valid_reg;
  reg  blockRefill_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
  wire  blockRefill_t = blockRefill ^ blockRefill_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
  wire  toggle_6582_clock;
  wire  toggle_6582_reset;
  wire  toggle_6582_valid;
  reg  toggle_6582_valid_reg;
  GEN_w64_toggle #(.COVER_INDEX(6197)) toggle_6197 (
    .clock(toggle_6197_clock),
    .reset(toggle_6197_reset),
    .valid(toggle_6197_valid)
  );
  GEN_w3_toggle #(.COVER_INDEX(6261)) toggle_6261 (
    .clock(toggle_6261_clock),
    .reset(toggle_6261_reset),
    .valid(toggle_6261_valid)
  );
  GEN_w2_toggle #(.COVER_INDEX(6264)) toggle_6264 (
    .clock(toggle_6264_clock),
    .reset(toggle_6264_reset),
    .valid(toggle_6264_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(6266)) toggle_6266 (
    .clock(toggle_6266_clock),
    .reset(toggle_6266_reset),
    .valid(toggle_6266_valid)
  );
  GEN_w18_toggle #(.COVER_INDEX(6330)) toggle_6330 (
    .clock(toggle_6330_clock),
    .reset(toggle_6330_reset),
    .valid(toggle_6330_valid)
  );
  GEN_w56_toggle #(.COVER_INDEX(6348)) toggle_6348 (
    .clock(toggle_6348_clock),
    .reset(toggle_6348_reset),
    .valid(toggle_6348_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(6404)) toggle_6404 (
    .clock(toggle_6404_clock),
    .reset(toggle_6404_reset),
    .valid(toggle_6404_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(6405)) toggle_6405 (
    .clock(toggle_6405_clock),
    .reset(toggle_6405_reset),
    .valid(toggle_6405_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(6406)) toggle_6406 (
    .clock(toggle_6406_clock),
    .reset(toggle_6406_reset),
    .valid(toggle_6406_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(6407)) toggle_6407 (
    .clock(toggle_6407_clock),
    .reset(toggle_6407_reset),
    .valid(toggle_6407_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(6408)) toggle_6408 (
    .clock(toggle_6408_clock),
    .reset(toggle_6408_reset),
    .valid(toggle_6408_valid)
  );
  GEN_w4_toggle #(.COVER_INDEX(6409)) toggle_6409 (
    .clock(toggle_6409_clock),
    .reset(toggle_6409_reset),
    .valid(toggle_6409_valid)
  );
  GEN_w27_toggle #(.COVER_INDEX(6413)) toggle_6413 (
    .clock(toggle_6413_clock),
    .reset(toggle_6413_reset),
    .valid(toggle_6413_valid)
  );
  GEN_w16_toggle #(.COVER_INDEX(6440)) toggle_6440 (
    .clock(toggle_6440_clock),
    .reset(toggle_6440_reset),
    .valid(toggle_6440_valid)
  );
  GEN_w18_toggle #(.COVER_INDEX(6456)) toggle_6456 (
    .clock(toggle_6456_clock),
    .reset(toggle_6456_reset),
    .valid(toggle_6456_valid)
  );
  GEN_w8_toggle #(.COVER_INDEX(6474)) toggle_6474 (
    .clock(toggle_6474_clock),
    .reset(toggle_6474_reset),
    .valid(toggle_6474_valid)
  );
  GEN_w44_toggle #(.COVER_INDEX(6482)) toggle_6482 (
    .clock(toggle_6482_clock),
    .reset(toggle_6482_reset),
    .valid(toggle_6482_valid)
  );
  GEN_w56_toggle #(.COVER_INDEX(6526)) toggle_6526 (
    .clock(toggle_6526_clock),
    .reset(toggle_6526_reset),
    .valid(toggle_6526_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(6582)) toggle_6582 (
    .clock(toggle_6582_clock),
    .reset(toggle_6582_reset),
    .valid(toggle_6582_valid)
  );
  assign io_in_ready = io_out_ready & _T_35 & ~miss & io_mdReady & _io_out_valid_T_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 498:86]
  assign io_out_valid = out_req_valid & ~hasException; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 496:75]
  assign io_out_bits_addr = paddr[31:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 483:20]
  assign io_out_bits_user = io_in_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 482:15]
  assign io_mdWrite_wen = blockRefill ? 1'h0 : REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 454:22 455:20 src/main/scala/nutcore/mem/TLB.scala 217:14]
  assign io_mdWrite_waymask = REG_2; // @[src/main/scala/nutcore/mem/TLB.scala 219:18]
  assign io_mdWrite_wdata = _io_mdWrite_wdata_T[144:0]; // @[src/main/scala/nutcore/mem/TLB.scala 220:16]
  assign io_mem_req_valid = (state == 3'h1 | cmd) & ~isFlush & ~raddrCancel; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 442:85]
  assign io_mem_req_bits_addr = raddr[31:0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_mem_req_bits_cmd = {{3'd0}, cmd}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 441:138]
  assign io_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 443:21]
  assign io_pf_loadPF = 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:16]
  assign io_pf_storePF = 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 285:17]
  assign io_pf_laf = 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:13]
  assign io_pf_saf = 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:13]
  assign io_ipf = hit ? hitinstrPF : missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 500:16]
  assign io_iaf = out_req_valid & (~_instrAF_T_7 | missPTEAF); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 486:30]
  assign io_isFinish = _alreadyOutFire_T | hasException; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 502:32]
  assign toggle_6197_clock = clock;
  assign toggle_6197_reset = reset;
  assign toggle_6197_valid = victimWaymask_lfsr ^ toggle_6197_valid_reg;
  assign toggle_6261_clock = clock;
  assign toggle_6261_reset = reset;
  assign toggle_6261_valid = state ^ toggle_6261_valid_reg;
  assign toggle_6264_clock = clock;
  assign toggle_6264_reset = reset;
  assign toggle_6264_valid = level ^ toggle_6264_valid_reg;
  assign toggle_6266_clock = clock;
  assign toggle_6266_reset = reset;
  assign toggle_6266_valid = memRespStore ^ toggle_6266_valid_reg;
  assign toggle_6330_clock = clock;
  assign toggle_6330_reset = reset;
  assign toggle_6330_valid = missMaskStore ^ toggle_6330_valid_reg;
  assign toggle_6348_clock = clock;
  assign toggle_6348_reset = reset;
  assign toggle_6348_valid = raddr ^ toggle_6348_valid_reg;
  assign toggle_6404_clock = clock;
  assign toggle_6404_reset = reset;
  assign toggle_6404_valid = alreadyOutFire ^ toggle_6404_valid_reg;
  assign toggle_6405_clock = clock;
  assign toggle_6405_reset = reset;
  assign toggle_6405_valid = needFlush ^ toggle_6405_valid_reg;
  assign toggle_6406_clock = clock;
  assign toggle_6406_reset = reset;
  assign toggle_6406_valid = missIPF ^ toggle_6406_valid_reg;
  assign toggle_6407_clock = clock;
  assign toggle_6407_reset = reset;
  assign toggle_6407_valid = missPTEAF ^ toggle_6407_valid_reg;
  assign toggle_6408_clock = clock;
  assign toggle_6408_reset = reset;
  assign toggle_6408_valid = REG ^ toggle_6408_valid_reg;
  assign toggle_6409_clock = clock;
  assign toggle_6409_reset = reset;
  assign toggle_6409_valid = REG_2 ^ toggle_6409_valid_reg;
  assign toggle_6413_clock = clock;
  assign toggle_6413_reset = reset;
  assign toggle_6413_valid = REG_3 ^ toggle_6413_valid_reg;
  assign toggle_6440_clock = clock;
  assign toggle_6440_reset = reset;
  assign toggle_6440_valid = REG_4 ^ toggle_6440_valid_reg;
  assign toggle_6456_clock = clock;
  assign toggle_6456_reset = reset;
  assign toggle_6456_valid = REG_5 ^ toggle_6456_valid_reg;
  assign toggle_6474_clock = clock;
  assign toggle_6474_reset = reset;
  assign toggle_6474_valid = REG_6 ^ toggle_6474_valid_reg;
  assign toggle_6482_clock = clock;
  assign toggle_6482_reset = reset;
  assign toggle_6482_valid = REG_7 ^ toggle_6482_valid_reg;
  assign toggle_6526_clock = clock;
  assign toggle_6526_reset = reset;
  assign toggle_6526_valid = REG_8 ^ toggle_6526_valid_reg;
  assign toggle_6582_clock = clock;
  assign toggle_6582_reset = reset;
  assign toggle_6582_valid = blockRefill ^ toggle_6582_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/LFSR64.scala 25:23]
      victimWaymask_lfsr <= 64'h1234567887654321; // @[src/main/scala/utils/LFSR64.scala 25:23]
    end else if (victimWaymask_lfsr == 64'h0) begin // @[src/main/scala/utils/LFSR64.scala 28:18]
      victimWaymask_lfsr <= 64'h1;
    end else begin
      victimWaymask_lfsr <= _victimWaymask_lfsr_T_2;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
      state <= 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        state <= 3'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 329:15]
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (isFlush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 338:22]
        state <= 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 339:15]
      end else begin
        state <= _GEN_17;
      end
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      state <= _GEN_53;
    end else begin
      state <= _GEN_75;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
      level <= 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        level <= 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 331:15]
      end
    end else if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        level <= _GEN_62;
      end
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
          if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
            memRespStore <= _GEN_49;
          end
        end
      end
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
          if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
            missMaskStore <= _GEN_52;
          end
        end
      end
    end
    if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        raddr <= _raddr_T_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 330:15]
      end
    end else if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
          raddr <= _GEN_47;
        end
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 333:24]
      end else begin
        alreadyOutFire <= _GEN_2;
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      alreadyOutFire <= _GEN_2;
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      alreadyOutFire <= _GEN_2;
    end else begin
      alreadyOutFire <= _GEN_79;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 312:26]
      needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 312:26]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss & _T_5) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 332:19]
      end else begin
        needFlush <= _GEN_4;
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (isFlush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 338:22]
        needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 340:19]
      end else begin
        needFlush <= _GEN_4;
      end
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      needFlush <= _GEN_54;
    end else begin
      needFlush <= _GEN_76;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24]
      missIPF <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24]
    end else if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
          missIPF <= _GEN_55;
        end else begin
          missIPF <= _GEN_77;
        end
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
      missPTEAF <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
    end else if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (!(isFlush)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 338:22]
          missPTEAF <= _GEN_18;
        end
      end else if (!(3'h2 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        missPTEAF <= _GEN_78;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
      REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
    end else begin
      REG <= missMetaRefill & _io_mem_req_valid_T_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
    end
    if (hit) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:20]
      REG_2 <= hitVec;
    end else begin
      REG_2 <= victimWaymask;
    end
    REG_3 <= {hitVec_hi,vpn_vpn0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:89]
    REG_4 <= io_satp[59:44]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 244:30]
    if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
        REG_5 <= _GEN_51;
      end else begin
        REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
      end
    end else begin
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
    end
    if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
        REG_6 <= _GEN_48;
      end else begin
        REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
      end
    end else begin
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
    end
    REG_7 <= io_mem_resp_bits_rdata[53:10]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
    REG_8 <= raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:27]
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
      blockRefill <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
    end else begin
      blockRefill <= _T_34 & mdMayHasAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    victimWaymask_lfsr_p <= victimWaymask_lfsr; // @[src/main/scala/utils/LFSR64.scala 25:23]
    toggle_6197_valid_reg <= victimWaymask_lfsr;
    state_p <= state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
    toggle_6261_valid_reg <= state;
    level_p <= level; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
    toggle_6264_valid_reg <= level;
    memRespStore_p <= memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    toggle_6266_valid_reg <= memRespStore;
    missMaskStore_p <= missMaskStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    toggle_6330_valid_reg <= missMaskStore;
    raddr_p <= raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    toggle_6348_valid_reg <= raddr;
    alreadyOutFire_p <= alreadyOutFire; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
    toggle_6404_valid_reg <= alreadyOutFire;
    needFlush_p <= needFlush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 312:26]
    toggle_6405_valid_reg <= needFlush;
    missIPF_p <= missIPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24]
    toggle_6406_valid_reg <= missIPF;
    missPTEAF_p <= missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
    toggle_6407_valid_reg <= missPTEAF;
    REG_p <= REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
    toggle_6408_valid_reg <= REG;
    REG_2_p <= REG_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:60]
    toggle_6409_valid_reg <= REG_2;
    REG_3_p <= REG_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    toggle_6413_valid_reg <= REG_3;
    REG_4_p <= REG_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    toggle_6440_valid_reg <= REG_4;
    REG_5_p <= REG_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    toggle_6456_valid_reg <= REG_5;
    REG_6_p <= REG_6; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
    toggle_6474_valid_reg <= REG_6;
    REG_7_p <= REG_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    toggle_6482_valid_reg <= REG_7;
    REG_8_p <= REG_8; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    toggle_6526_valid_reg <= REG_8;
    blockRefill_p <= blockRefill; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
    toggle_6582_valid_reg <= blockRefill;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  victimWaymask_lfsr = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  level = _RAND_2[1:0];
  _RAND_3 = {2{`RANDOM}};
  memRespStore = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  missMaskStore = _RAND_4[17:0];
  _RAND_5 = {2{`RANDOM}};
  raddr = _RAND_5[55:0];
  _RAND_6 = {1{`RANDOM}};
  alreadyOutFire = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  needFlush = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  missIPF = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  missPTEAF = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  REG = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  REG_2 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  REG_3 = _RAND_12[26:0];
  _RAND_13 = {1{`RANDOM}};
  REG_4 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  REG_5 = _RAND_14[17:0];
  _RAND_15 = {1{`RANDOM}};
  REG_6 = _RAND_15[7:0];
  _RAND_16 = {2{`RANDOM}};
  REG_7 = _RAND_16[43:0];
  _RAND_17 = {2{`RANDOM}};
  REG_8 = _RAND_17[55:0];
  _RAND_18 = {1{`RANDOM}};
  blockRefill = _RAND_18[0:0];
  _RAND_19 = {2{`RANDOM}};
  victimWaymask_lfsr_p = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  toggle_6197_valid_reg = _RAND_20[63:0];
  _RAND_21 = {1{`RANDOM}};
  state_p = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  toggle_6261_valid_reg = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  level_p = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  toggle_6264_valid_reg = _RAND_24[1:0];
  _RAND_25 = {2{`RANDOM}};
  memRespStore_p = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  toggle_6266_valid_reg = _RAND_26[63:0];
  _RAND_27 = {1{`RANDOM}};
  missMaskStore_p = _RAND_27[17:0];
  _RAND_28 = {1{`RANDOM}};
  toggle_6330_valid_reg = _RAND_28[17:0];
  _RAND_29 = {2{`RANDOM}};
  raddr_p = _RAND_29[55:0];
  _RAND_30 = {2{`RANDOM}};
  toggle_6348_valid_reg = _RAND_30[55:0];
  _RAND_31 = {1{`RANDOM}};
  alreadyOutFire_p = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  toggle_6404_valid_reg = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  needFlush_p = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  toggle_6405_valid_reg = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  missIPF_p = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  toggle_6406_valid_reg = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  missPTEAF_p = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  toggle_6407_valid_reg = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  REG_p = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  toggle_6408_valid_reg = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  REG_2_p = _RAND_41[3:0];
  _RAND_42 = {1{`RANDOM}};
  toggle_6409_valid_reg = _RAND_42[3:0];
  _RAND_43 = {1{`RANDOM}};
  REG_3_p = _RAND_43[26:0];
  _RAND_44 = {1{`RANDOM}};
  toggle_6413_valid_reg = _RAND_44[26:0];
  _RAND_45 = {1{`RANDOM}};
  REG_4_p = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  toggle_6440_valid_reg = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  REG_5_p = _RAND_47[17:0];
  _RAND_48 = {1{`RANDOM}};
  toggle_6456_valid_reg = _RAND_48[17:0];
  _RAND_49 = {1{`RANDOM}};
  REG_6_p = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  toggle_6474_valid_reg = _RAND_50[7:0];
  _RAND_51 = {2{`RANDOM}};
  REG_7_p = _RAND_51[43:0];
  _RAND_52 = {2{`RANDOM}};
  toggle_6482_valid_reg = _RAND_52[43:0];
  _RAND_53 = {2{`RANDOM}};
  REG_8_p = _RAND_53[55:0];
  _RAND_54 = {2{`RANDOM}};
  toggle_6526_valid_reg = _RAND_54[55:0];
  _RAND_55 = {1{`RANDOM}};
  blockRefill_p = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  toggle_6582_valid_reg = _RAND_56[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[0]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[1]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[2]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[3]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[4]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[5]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[6]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[7]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[8]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[9]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[10]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[11]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[12]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[13]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[14]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[15]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[16]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[17]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[18]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[19]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[20]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[21]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[22]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[23]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[24]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[25]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[26]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[27]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[28]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[29]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[30]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[31]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[32]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[33]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[34]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[35]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[36]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[37]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[38]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[39]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[40]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[41]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[42]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[43]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[44]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[45]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[46]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[47]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[48]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[49]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[50]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[51]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[52]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[53]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[54]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[55]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[56]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[57]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[58]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[59]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[60]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[61]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[62]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[63]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(state_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
    end
    //
    if (enToggle_past) begin
      cover(level_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
    end
    //
    if (enToggle_past) begin
      cover(level_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[39]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[40]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[41]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[42]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[43]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[44]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[45]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[46]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[47]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[48]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[49]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[50]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[51]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[52]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[53]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[54]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[55]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[56]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[57]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[58]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[59]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[60]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[61]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[62]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[63]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[39]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[40]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[41]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[42]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[43]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[44]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[45]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[46]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[47]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[48]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[49]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[50]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[51]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[52]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[53]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[54]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[55]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(alreadyOutFire_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
    end
    //
    if (enToggle_past) begin
      cover(needFlush_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 312:26]
    end
    //
    if (enToggle_past) begin
      cover(missIPF_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 318:24]
    end
    //
    if (enToggle_past) begin
      cover(missPTEAF_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(REG_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
    end
    //
    if (enToggle_past) begin
      cover(REG_2_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:60]
    end
    //
    if (enToggle_past) begin
      cover(REG_2_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:60]
    end
    //
    if (enToggle_past) begin
      cover(REG_2_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:60]
    end
    //
    if (enToggle_past) begin
      cover(REG_2_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:60]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_6_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_6_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_6_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_6_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_6_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_6_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_6_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_6_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[39]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[40]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[41]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[42]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[43]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[39]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[40]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[41]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[42]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[43]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[44]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[45]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[46]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[47]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[48]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[49]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[50]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[51]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[52]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[53]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[54]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[55]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(blockRefill_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
    end
  end
endmodule
module EmbeddedTLBEmpty(
  input   clock,
  input   reset
);
endmodule
module EmbeddedTLBMD(
  input          clock,
  input          reset,
  output [144:0] io_tlbmd_0, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output [144:0] io_tlbmd_1, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output [144:0] io_tlbmd_2, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output [144:0] io_tlbmd_3, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input          io_write_wen, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input  [3:0]   io_write_waymask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input  [144:0] io_write_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output         io_ready // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [159:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [144:0] tlbmd_0 [0:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_0_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_0_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg [144:0] tlbmd_1 [0:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_1_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_1_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg [144:0] tlbmd_2 [0:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_2_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_2_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg [144:0] tlbmd_3 [0:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_3_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_3_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg  resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 56:27]
  wire  _GEN_1 = resetState ? 1'h0 : resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 58:22 56:27 58:35]
  wire [3:0] waymask = resetState ? 4'hf : io_write_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 67:20]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  resetState_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 56:27]
  wire  resetState_t = resetState ^ resetState_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 56:27]
  wire  toggle_6583_clock;
  wire  toggle_6583_reset;
  wire  toggle_6583_valid;
  reg  toggle_6583_valid_reg;
  GEN_w1_toggle #(.COVER_INDEX(6583)) toggle_6583 (
    .clock(toggle_6583_clock),
    .reset(toggle_6583_reset),
    .valid(toggle_6583_valid)
  );
  assign tlbmd_0_MPORT_en = 1'h1;
  assign tlbmd_0_MPORT_addr = 1'h0;
  assign tlbmd_0_MPORT_data = tlbmd_0[tlbmd_0_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_0_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_0_MPORT_1_addr = 1'h0;
  assign tlbmd_0_MPORT_1_mask = waymask[0];
  assign tlbmd_0_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_1_MPORT_en = 1'h1;
  assign tlbmd_1_MPORT_addr = 1'h0;
  assign tlbmd_1_MPORT_data = tlbmd_1[tlbmd_1_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_1_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_1_MPORT_1_addr = 1'h0;
  assign tlbmd_1_MPORT_1_mask = waymask[1];
  assign tlbmd_1_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_2_MPORT_en = 1'h1;
  assign tlbmd_2_MPORT_addr = 1'h0;
  assign tlbmd_2_MPORT_data = tlbmd_2[tlbmd_2_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_2_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_2_MPORT_1_addr = 1'h0;
  assign tlbmd_2_MPORT_1_mask = waymask[2];
  assign tlbmd_2_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_3_MPORT_en = 1'h1;
  assign tlbmd_3_MPORT_addr = 1'h0;
  assign tlbmd_3_MPORT_data = tlbmd_3[tlbmd_3_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_3_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_3_MPORT_1_addr = 1'h0;
  assign tlbmd_3_MPORT_1_mask = waymask[3];
  assign tlbmd_3_MPORT_1_en = resetState | io_write_wen;
  assign io_tlbmd_0 = tlbmd_0_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_tlbmd_1 = tlbmd_1_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_tlbmd_2 = tlbmd_2_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_tlbmd_3 = tlbmd_3_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_ready = ~resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 73:15]
  assign toggle_6583_clock = clock;
  assign toggle_6583_reset = reset;
  assign toggle_6583_valid = resetState ^ toggle_6583_valid_reg;
  always @(posedge clock) begin
    if (tlbmd_0_MPORT_1_en & tlbmd_0_MPORT_1_mask) begin
      tlbmd_0[tlbmd_0_MPORT_1_addr] <= tlbmd_0_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    if (tlbmd_1_MPORT_1_en & tlbmd_1_MPORT_1_mask) begin
      tlbmd_1[tlbmd_1_MPORT_1_addr] <= tlbmd_1_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    if (tlbmd_2_MPORT_1_en & tlbmd_2_MPORT_1_mask) begin
      tlbmd_2[tlbmd_2_MPORT_1_addr] <= tlbmd_2_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    if (tlbmd_3_MPORT_1_en & tlbmd_3_MPORT_1_mask) begin
      tlbmd_3[tlbmd_3_MPORT_1_addr] <= tlbmd_3_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    resetState <= reset | _GEN_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 56:{27,27}]
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    resetState_p <= resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 56:27]
    toggle_6583_valid_reg <= resetState;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {5{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_0[initvar] = _RAND_0[144:0];
  _RAND_1 = {5{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_1[initvar] = _RAND_1[144:0];
  _RAND_2 = {5{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_2[initvar] = _RAND_2[144:0];
  _RAND_3 = {5{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_3[initvar] = _RAND_3[144:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  resetState = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  resetState_p = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  toggle_6583_valid_reg = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(resetState_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 56:27]
    end
  end
endmodule
module EmbeddedTLB(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [38:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [86:0] io_in_req_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_in_resp_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [86:0] io_in_resp_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_out_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_out_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [86:0] io_out_req_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_out_resp_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_out_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [63:0] io_out_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [86:0] io_out_resp_bits_user, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_mem_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_mem_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [31:0] io_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [3:0]  io_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [63:0] io_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_mem_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [63:0] io_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_flush, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [1:0]  io_csrMMU_priviledgeMode, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_iaf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [63:0] CSRSATP,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [159:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [95:0] _RAND_9;
  reg [95:0] _RAND_10;
  reg [159:0] _RAND_11;
  reg [159:0] _RAND_12;
  reg [159:0] _RAND_13;
  reg [159:0] _RAND_14;
  reg [159:0] _RAND_15;
  reg [159:0] _RAND_16;
  reg [159:0] _RAND_17;
  reg [159:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [95:0] _RAND_29;
  reg [95:0] _RAND_30;
  reg [95:0] _RAND_31;
  reg [95:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  wire  tlbExec_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_in_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [38:0] tlbExec_io_in_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [86:0] tlbExec_io_in_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_out_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_out_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [31:0] tlbExec_io_out_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [86:0] tlbExec_io_out_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mdWrite_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_mdWrite_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_mdWrite_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mdReady; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [31:0] tlbExec_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_satp; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [1:0] tlbExec_io_pf_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_laf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_saf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_ipf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_iaf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_isFinish; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbEmpty_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire  tlbEmpty_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire  mdTLB_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  mdTLB_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  mdTLB_io_write_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [3:0] mdTLB_io_write_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_write_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  mdTLB_io_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  vmEnable = CSRSATP[63:60] == 4'h8 & io_csrMMU_priviledgeMode < 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 90:57]
  reg [144:0] r_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  reg [144:0] r_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  reg [144:0] r_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  reg [144:0] r_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire  mdUpdate = io_in_req_valid & tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:26]
  wire  _reqIsLegalInstr_T_2 = io_in_req_bits_addr >= 39'h40000000 & io_in_req_bits_addr < 39'h40001000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _reqIsLegalInstr_T_5 = io_in_req_bits_addr >= 39'h80000000 & io_in_req_bits_addr < 39'h100000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [1:0] _reqIsLegalInstr_T_6 = {_reqIsLegalInstr_T_5,_reqIsLegalInstr_T_2}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _reqIsLegalInstr_T_7 = |_reqIsLegalInstr_T_6; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  reqIsLegalInstr = vmEnable | _reqIsLegalInstr_T_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 119:34]
  reg  hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 120:28]
  wire  _lastReqAddr_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _lastReqAddr_T_2 = _lastReqAddr_T & ~io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:67]
  reg [38:0] lastReqAddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
  wire  _T_1 = io_in_resp_ready & io_in_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _GEN_5 = _T_1 & io_in_resp_bits_user[38:0] == lastReqAddr ? 1'h0 : hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 127:96 128:19 120:28]
  wire  _GEN_6 = _lastReqAddr_T | _GEN_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 125:33 126:19]
  reg  hasIllegalInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 131:35]
  wire  _hasIllegalInflight_T = ~reqIsLegalInstr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 135:27]
  reg  valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
  wire  _GEN_10 = tlbExec_io_isFinish ? 1'h0 : valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24 108:{25,33}]
  wire  _GEN_11 = mdUpdate & vmEnable | _GEN_10; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 109:{50,58}]
  reg [38:0] tlbExec_io_in_bits_r_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  reg [86:0] tlbExec_io_in_bits_r_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  wire  _GEN_19 = io_in_req_valid & _hasIllegalInflight_T ? ~hasInflight : io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 157:23 158:50 159:25]
  wire  _GEN_20 = ~vmEnable | io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 145:26 170:23]
  wire  _GEN_21 = ~vmEnable ? io_in_req_valid & reqIsLegalInstr : tlbExec_io_out_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 156:24 170:23]
  reg [86:0] userBits; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [144:0] r_0_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire [144:0] r_0_t = r_0 ^ r_0_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire  toggle_6584_clock;
  wire  toggle_6584_reset;
  wire [144:0] toggle_6584_valid;
  reg [144:0] toggle_6584_valid_reg;
  reg [144:0] r_1_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire [144:0] r_1_t = r_1 ^ r_1_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire  toggle_6729_clock;
  wire  toggle_6729_reset;
  wire [144:0] toggle_6729_valid;
  reg [144:0] toggle_6729_valid_reg;
  reg [144:0] r_2_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire [144:0] r_2_t = r_2 ^ r_2_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire  toggle_6874_clock;
  wire  toggle_6874_reset;
  wire [144:0] toggle_6874_valid;
  reg [144:0] toggle_6874_valid_reg;
  reg [144:0] r_3_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire [144:0] r_3_t = r_3 ^ r_3_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire  toggle_7019_clock;
  wire  toggle_7019_reset;
  wire [144:0] toggle_7019_valid;
  reg [144:0] toggle_7019_valid_reg;
  reg  hasInflight_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 120:28]
  wire  hasInflight_t = hasInflight ^ hasInflight_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 120:28]
  wire  toggle_7164_clock;
  wire  toggle_7164_reset;
  wire  toggle_7164_valid;
  reg  toggle_7164_valid_reg;
  reg [38:0] lastReqAddr_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
  wire [38:0] lastReqAddr_t = lastReqAddr ^ lastReqAddr_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
  wire  toggle_7165_clock;
  wire  toggle_7165_reset;
  wire [38:0] toggle_7165_valid;
  reg [38:0] toggle_7165_valid_reg;
  reg  hasIllegalInflight_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 131:35]
  wire  hasIllegalInflight_t = hasIllegalInflight ^ hasIllegalInflight_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 131:35]
  wire  toggle_7204_clock;
  wire  toggle_7204_reset;
  wire  toggle_7204_valid;
  reg  toggle_7204_valid_reg;
  reg  valid_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
  wire  valid_t = valid ^ valid_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
  wire  toggle_7205_clock;
  wire  toggle_7205_reset;
  wire  toggle_7205_valid;
  reg  toggle_7205_valid_reg;
  reg [38:0] tlbExec_io_in_bits_r_addr_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  wire [38:0] tlbExec_io_in_bits_r_addr_t = tlbExec_io_in_bits_r_addr ^ tlbExec_io_in_bits_r_addr_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  wire  toggle_7206_clock;
  wire  toggle_7206_reset;
  wire [38:0] toggle_7206_valid;
  reg [38:0] toggle_7206_valid_reg;
  reg [86:0] tlbExec_io_in_bits_r_user_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  wire [86:0] tlbExec_io_in_bits_r_user_t = tlbExec_io_in_bits_r_user ^ tlbExec_io_in_bits_r_user_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  wire  toggle_7245_clock;
  wire  toggle_7245_reset;
  wire [86:0] toggle_7245_valid;
  reg [86:0] toggle_7245_valid_reg;
  reg [86:0] userBits_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
  wire [86:0] userBits_t = userBits ^ userBits_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
  wire  toggle_7332_clock;
  wire  toggle_7332_reset;
  wire [86:0] toggle_7332_valid;
  reg [86:0] toggle_7332_valid_reg;
  EmbeddedTLBExec tlbExec ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
    .clock(tlbExec_clock),
    .reset(tlbExec_reset),
    .io_in_ready(tlbExec_io_in_ready),
    .io_in_valid(tlbExec_io_in_valid),
    .io_in_bits_addr(tlbExec_io_in_bits_addr),
    .io_in_bits_user(tlbExec_io_in_bits_user),
    .io_out_ready(tlbExec_io_out_ready),
    .io_out_valid(tlbExec_io_out_valid),
    .io_out_bits_addr(tlbExec_io_out_bits_addr),
    .io_out_bits_user(tlbExec_io_out_bits_user),
    .io_md_0(tlbExec_io_md_0),
    .io_md_1(tlbExec_io_md_1),
    .io_md_2(tlbExec_io_md_2),
    .io_md_3(tlbExec_io_md_3),
    .io_mdWrite_wen(tlbExec_io_mdWrite_wen),
    .io_mdWrite_waymask(tlbExec_io_mdWrite_waymask),
    .io_mdWrite_wdata(tlbExec_io_mdWrite_wdata),
    .io_mdReady(tlbExec_io_mdReady),
    .io_mem_req_ready(tlbExec_io_mem_req_ready),
    .io_mem_req_valid(tlbExec_io_mem_req_valid),
    .io_mem_req_bits_addr(tlbExec_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(tlbExec_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(tlbExec_io_mem_req_bits_wdata),
    .io_mem_resp_ready(tlbExec_io_mem_resp_ready),
    .io_mem_resp_valid(tlbExec_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(tlbExec_io_mem_resp_bits_rdata),
    .io_flush(tlbExec_io_flush),
    .io_satp(tlbExec_io_satp),
    .io_pf_priviledgeMode(tlbExec_io_pf_priviledgeMode),
    .io_pf_loadPF(tlbExec_io_pf_loadPF),
    .io_pf_storePF(tlbExec_io_pf_storePF),
    .io_pf_laf(tlbExec_io_pf_laf),
    .io_pf_saf(tlbExec_io_pf_saf),
    .io_ipf(tlbExec_io_ipf),
    .io_iaf(tlbExec_io_iaf),
    .io_isFinish(tlbExec_io_isFinish)
  );
  EmbeddedTLBEmpty tlbEmpty ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
    .clock(tlbEmpty_clock),
    .reset(tlbEmpty_reset)
  );
  EmbeddedTLBMD mdTLB ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
    .clock(mdTLB_clock),
    .reset(mdTLB_reset),
    .io_tlbmd_0(mdTLB_io_tlbmd_0),
    .io_tlbmd_1(mdTLB_io_tlbmd_1),
    .io_tlbmd_2(mdTLB_io_tlbmd_2),
    .io_tlbmd_3(mdTLB_io_tlbmd_3),
    .io_write_wen(mdTLB_io_write_wen),
    .io_write_waymask(mdTLB_io_write_waymask),
    .io_write_wdata(mdTLB_io_write_wdata),
    .io_ready(mdTLB_io_ready)
  );
  GEN_w145_toggle #(.COVER_INDEX(6584)) toggle_6584 (
    .clock(toggle_6584_clock),
    .reset(toggle_6584_reset),
    .valid(toggle_6584_valid)
  );
  GEN_w145_toggle #(.COVER_INDEX(6729)) toggle_6729 (
    .clock(toggle_6729_clock),
    .reset(toggle_6729_reset),
    .valid(toggle_6729_valid)
  );
  GEN_w145_toggle #(.COVER_INDEX(6874)) toggle_6874 (
    .clock(toggle_6874_clock),
    .reset(toggle_6874_reset),
    .valid(toggle_6874_valid)
  );
  GEN_w145_toggle #(.COVER_INDEX(7019)) toggle_7019 (
    .clock(toggle_7019_clock),
    .reset(toggle_7019_reset),
    .valid(toggle_7019_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(7164)) toggle_7164 (
    .clock(toggle_7164_clock),
    .reset(toggle_7164_reset),
    .valid(toggle_7164_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(7165)) toggle_7165 (
    .clock(toggle_7165_clock),
    .reset(toggle_7165_reset),
    .valid(toggle_7165_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(7204)) toggle_7204 (
    .clock(toggle_7204_clock),
    .reset(toggle_7204_reset),
    .valid(toggle_7204_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(7205)) toggle_7205 (
    .clock(toggle_7205_clock),
    .reset(toggle_7205_reset),
    .valid(toggle_7205_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(7206)) toggle_7206 (
    .clock(toggle_7206_clock),
    .reset(toggle_7206_reset),
    .valid(toggle_7206_valid)
  );
  GEN_w87_toggle #(.COVER_INDEX(7245)) toggle_7245 (
    .clock(toggle_7245_clock),
    .reset(toggle_7245_reset),
    .valid(toggle_7245_valid)
  );
  GEN_w87_toggle #(.COVER_INDEX(7332)) toggle_7332 (
    .clock(toggle_7332_clock),
    .reset(toggle_7332_reset),
    .valid(toggle_7332_valid)
  );
  assign io_in_req_ready = ~vmEnable ? _GEN_19 : tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 112:16 144:19]
  assign io_in_resp_valid = hasIllegalInflight & io_iaf | io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 201:41 202:24]
  assign io_in_resp_bits_rdata = hasIllegalInflight & io_iaf ? 64'h0 : io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 201:41 203:29]
  assign io_in_resp_bits_user = hasIllegalInflight & io_iaf ? userBits : io_out_resp_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 201:41 206:34]
  assign io_out_req_valid = (tlbExec_io_ipf | tlbExec_io_iaf) & vmEnable ? 1'h0 : _GEN_21; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 189:59 191:24]
  assign io_out_req_bits_addr = ~vmEnable ? io_in_req_bits_addr[31:0] : tlbExec_io_out_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 162:26 170:23]
  assign io_out_req_bits_user = ~vmEnable ? io_in_req_bits_user : tlbExec_io_out_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 167:32 170:23]
  assign io_out_resp_ready = io_in_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 172:15]
  assign io_mem_req_valid = tlbExec_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_mem_req_bits_addr = tlbExec_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_mem_req_bits_cmd = tlbExec_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_mem_req_bits_wdata = tlbExec_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_iaf = vmEnable ? tlbExec_io_iaf : hasIllegalInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 212:16]
  assign tlbExec_clock = clock;
  assign tlbExec_reset = reset;
  assign tlbExec_io_in_valid = valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 114:17]
  assign tlbExec_io_in_bits_addr = tlbExec_io_in_bits_r_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_in_bits_user = tlbExec_io_in_bits_r_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_out_ready = (tlbExec_io_ipf | tlbExec_io_iaf) & vmEnable ? 1'h0 : _GEN_20; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 189:59 190:28]
  assign tlbExec_io_md_0 = r_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_md_1 = r_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_md_2 = r_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_md_3 = r_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_mdReady = mdTLB_io_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 97:22]
  assign tlbExec_io_mem_req_ready = io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign tlbExec_io_mem_resp_valid = io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign tlbExec_io_mem_resp_bits_rdata = io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign tlbExec_io_flush = io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 92:20]
  assign tlbExec_io_satp = CSRSATP; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 80:22]
  assign tlbExec_io_pf_priviledgeMode = io_csrMMU_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 95:17]
  assign tlbEmpty_clock = clock;
  assign tlbEmpty_reset = reset;
  assign mdTLB_clock = clock;
  assign mdTLB_reset = reset | MOUFlushTLB; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 104:31]
  assign mdTLB_io_write_wen = tlbExec_io_mdWrite_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  assign mdTLB_io_write_waymask = tlbExec_io_mdWrite_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  assign mdTLB_io_write_wdata = tlbExec_io_mdWrite_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  assign toggle_6584_clock = clock;
  assign toggle_6584_reset = reset;
  assign toggle_6584_valid = r_0 ^ toggle_6584_valid_reg;
  assign toggle_6729_clock = clock;
  assign toggle_6729_reset = reset;
  assign toggle_6729_valid = r_1 ^ toggle_6729_valid_reg;
  assign toggle_6874_clock = clock;
  assign toggle_6874_reset = reset;
  assign toggle_6874_valid = r_2 ^ toggle_6874_valid_reg;
  assign toggle_7019_clock = clock;
  assign toggle_7019_reset = reset;
  assign toggle_7019_valid = r_3 ^ toggle_7019_valid_reg;
  assign toggle_7164_clock = clock;
  assign toggle_7164_reset = reset;
  assign toggle_7164_valid = hasInflight ^ toggle_7164_valid_reg;
  assign toggle_7165_clock = clock;
  assign toggle_7165_reset = reset;
  assign toggle_7165_valid = lastReqAddr ^ toggle_7165_valid_reg;
  assign toggle_7204_clock = clock;
  assign toggle_7204_reset = reset;
  assign toggle_7204_valid = hasIllegalInflight ^ toggle_7204_valid_reg;
  assign toggle_7205_clock = clock;
  assign toggle_7205_reset = reset;
  assign toggle_7205_valid = valid ^ toggle_7205_valid_reg;
  assign toggle_7206_clock = clock;
  assign toggle_7206_reset = reset;
  assign toggle_7206_valid = tlbExec_io_in_bits_r_addr ^ toggle_7206_valid_reg;
  assign toggle_7245_clock = clock;
  assign toggle_7245_reset = reset;
  assign toggle_7245_valid = tlbExec_io_in_bits_r_user ^ toggle_7245_valid_reg;
  assign toggle_7332_clock = clock;
  assign toggle_7332_reset = reset;
  assign toggle_7332_valid = userBits ^ toggle_7332_valid_reg;
  always @(posedge clock) begin
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_0 <= mdTLB_io_tlbmd_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_1 <= mdTLB_io_tlbmd_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_2 <= mdTLB_io_tlbmd_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_3 <= mdTLB_io_tlbmd_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 120:28]
      hasInflight <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 120:28]
    end else if (io_flush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 123:21]
      hasInflight <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 124:19]
    end else begin
      hasInflight <= _GEN_6;
    end
    if (_lastReqAddr_T & ~io_flush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
      lastReqAddr <= io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 131:35]
      hasIllegalInflight <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 131:35]
    end else if (_T_1 | io_flush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 132:38]
      hasIllegalInflight <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 133:24]
    end else if (_lastReqAddr_T_2) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 134:44]
      hasIllegalInflight <= ~reqIsLegalInstr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 135:24]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
      valid <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
    end else if (io_flush) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 110:20]
      valid <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 110:28]
    end else begin
      valid <= _GEN_11;
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_addr <= io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_user <= io_in_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    if (_lastReqAddr_T_2) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
      userBits <= io_in_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    r_0_p <= r_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    toggle_6584_valid_reg <= r_0;
    r_1_p <= r_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    toggle_6729_valid_reg <= r_1;
    r_2_p <= r_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    toggle_6874_valid_reg <= r_2;
    r_3_p <= r_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    toggle_7019_valid_reg <= r_3;
    hasInflight_p <= hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 120:28]
    toggle_7164_valid_reg <= hasInflight;
    lastReqAddr_p <= lastReqAddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    toggle_7165_valid_reg <= lastReqAddr;
    hasIllegalInflight_p <= hasIllegalInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 131:35]
    toggle_7204_valid_reg <= hasIllegalInflight;
    valid_p <= valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
    toggle_7205_valid_reg <= valid;
    tlbExec_io_in_bits_r_addr_p <= tlbExec_io_in_bits_r_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    toggle_7206_valid_reg <= tlbExec_io_in_bits_r_addr;
    tlbExec_io_in_bits_r_user_p <= tlbExec_io_in_bits_r_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    toggle_7245_valid_reg <= tlbExec_io_in_bits_r_user;
    userBits_p <= userBits; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    toggle_7332_valid_reg <= userBits;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {5{`RANDOM}};
  r_0 = _RAND_0[144:0];
  _RAND_1 = {5{`RANDOM}};
  r_1 = _RAND_1[144:0];
  _RAND_2 = {5{`RANDOM}};
  r_2 = _RAND_2[144:0];
  _RAND_3 = {5{`RANDOM}};
  r_3 = _RAND_3[144:0];
  _RAND_4 = {1{`RANDOM}};
  hasInflight = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  lastReqAddr = _RAND_5[38:0];
  _RAND_6 = {1{`RANDOM}};
  hasIllegalInflight = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  valid = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  tlbExec_io_in_bits_r_addr = _RAND_8[38:0];
  _RAND_9 = {3{`RANDOM}};
  tlbExec_io_in_bits_r_user = _RAND_9[86:0];
  _RAND_10 = {3{`RANDOM}};
  userBits = _RAND_10[86:0];
  _RAND_11 = {5{`RANDOM}};
  r_0_p = _RAND_11[144:0];
  _RAND_12 = {5{`RANDOM}};
  toggle_6584_valid_reg = _RAND_12[144:0];
  _RAND_13 = {5{`RANDOM}};
  r_1_p = _RAND_13[144:0];
  _RAND_14 = {5{`RANDOM}};
  toggle_6729_valid_reg = _RAND_14[144:0];
  _RAND_15 = {5{`RANDOM}};
  r_2_p = _RAND_15[144:0];
  _RAND_16 = {5{`RANDOM}};
  toggle_6874_valid_reg = _RAND_16[144:0];
  _RAND_17 = {5{`RANDOM}};
  r_3_p = _RAND_17[144:0];
  _RAND_18 = {5{`RANDOM}};
  toggle_7019_valid_reg = _RAND_18[144:0];
  _RAND_19 = {1{`RANDOM}};
  hasInflight_p = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  toggle_7164_valid_reg = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  lastReqAddr_p = _RAND_21[38:0];
  _RAND_22 = {2{`RANDOM}};
  toggle_7165_valid_reg = _RAND_22[38:0];
  _RAND_23 = {1{`RANDOM}};
  hasIllegalInflight_p = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  toggle_7204_valid_reg = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  valid_p = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  toggle_7205_valid_reg = _RAND_26[0:0];
  _RAND_27 = {2{`RANDOM}};
  tlbExec_io_in_bits_r_addr_p = _RAND_27[38:0];
  _RAND_28 = {2{`RANDOM}};
  toggle_7206_valid_reg = _RAND_28[38:0];
  _RAND_29 = {3{`RANDOM}};
  tlbExec_io_in_bits_r_user_p = _RAND_29[86:0];
  _RAND_30 = {3{`RANDOM}};
  toggle_7245_valid_reg = _RAND_30[86:0];
  _RAND_31 = {3{`RANDOM}};
  userBits_p = _RAND_31[86:0];
  _RAND_32 = {3{`RANDOM}};
  toggle_7332_valid_reg = _RAND_32[86:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(r_0_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[39]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[40]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[41]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[42]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[43]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[44]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[45]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[46]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[47]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[48]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[49]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[50]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[51]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[52]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[53]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[54]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[55]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[56]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[57]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[58]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[59]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[60]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[61]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[62]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[63]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[64]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[65]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[66]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[67]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[68]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[69]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[70]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[71]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[72]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[73]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[74]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[75]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[76]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[77]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[78]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[79]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[80]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[81]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[82]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[83]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[84]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[85]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[86]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[87]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[88]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[89]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[90]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[91]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[92]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[93]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[94]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[95]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[96]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[97]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[98]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[99]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[100]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[101]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[102]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[103]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[104]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[105]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[106]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[107]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[108]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[109]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[110]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[111]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[112]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[113]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[114]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[115]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[116]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[117]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[118]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[119]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[120]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[121]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[122]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[123]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[124]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[125]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[126]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[127]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[128]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[129]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[130]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[131]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[132]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[133]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[134]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[135]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[136]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[137]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[138]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[139]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[140]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[141]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[142]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[143]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[144]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[39]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[40]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[41]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[42]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[43]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[44]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[45]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[46]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[47]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[48]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[49]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[50]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[51]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[52]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[53]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[54]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[55]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[56]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[57]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[58]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[59]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[60]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[61]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[62]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[63]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[64]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[65]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[66]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[67]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[68]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[69]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[70]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[71]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[72]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[73]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[74]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[75]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[76]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[77]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[78]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[79]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[80]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[81]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[82]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[83]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[84]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[85]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[86]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[87]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[88]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[89]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[90]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[91]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[92]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[93]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[94]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[95]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[96]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[97]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[98]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[99]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[100]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[101]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[102]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[103]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[104]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[105]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[106]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[107]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[108]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[109]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[110]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[111]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[112]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[113]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[114]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[115]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[116]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[117]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[118]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[119]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[120]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[121]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[122]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[123]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[124]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[125]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[126]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[127]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[128]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[129]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[130]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[131]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[132]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[133]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[134]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[135]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[136]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[137]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[138]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[139]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[140]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[141]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[142]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[143]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[144]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[39]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[40]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[41]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[42]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[43]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[44]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[45]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[46]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[47]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[48]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[49]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[50]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[51]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[52]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[53]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[54]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[55]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[56]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[57]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[58]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[59]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[60]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[61]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[62]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[63]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[64]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[65]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[66]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[67]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[68]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[69]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[70]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[71]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[72]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[73]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[74]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[75]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[76]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[77]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[78]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[79]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[80]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[81]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[82]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[83]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[84]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[85]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[86]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[87]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[88]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[89]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[90]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[91]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[92]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[93]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[94]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[95]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[96]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[97]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[98]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[99]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[100]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[101]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[102]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[103]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[104]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[105]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[106]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[107]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[108]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[109]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[110]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[111]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[112]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[113]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[114]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[115]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[116]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[117]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[118]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[119]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[120]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[121]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[122]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[123]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[124]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[125]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[126]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[127]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[128]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[129]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[130]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[131]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[132]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[133]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[134]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[135]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[136]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[137]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[138]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[139]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[140]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[141]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[142]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[143]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[144]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[39]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[40]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[41]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[42]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[43]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[44]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[45]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[46]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[47]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[48]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[49]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[50]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[51]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[52]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[53]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[54]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[55]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[56]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[57]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[58]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[59]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[60]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[61]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[62]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[63]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[64]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[65]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[66]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[67]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[68]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[69]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[70]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[71]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[72]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[73]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[74]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[75]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[76]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[77]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[78]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[79]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[80]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[81]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[82]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[83]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[84]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[85]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[86]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[87]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[88]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[89]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[90]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[91]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[92]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[93]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[94]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[95]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[96]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[97]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[98]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[99]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[100]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[101]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[102]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[103]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[104]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[105]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[106]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[107]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[108]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[109]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[110]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[111]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[112]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[113]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[114]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[115]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[116]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[117]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[118]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[119]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[120]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[121]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[122]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[123]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[124]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[125]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[126]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[127]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[128]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[129]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[130]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[131]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[132]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[133]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[134]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[135]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[136]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[137]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[138]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[139]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[140]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[141]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[142]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[143]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[144]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(hasInflight_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 120:28]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(lastReqAddr_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 121:30]
    end
    //
    if (enToggle_past) begin
      cover(hasIllegalInflight_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 131:35]
    end
    //
    if (enToggle_past) begin
      cover(valid_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[39]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[40]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[41]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[42]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[43]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[44]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[45]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[46]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[47]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[48]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[49]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[50]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[51]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[52]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[53]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[54]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[55]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[56]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[57]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[58]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[59]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[60]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[61]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[62]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[63]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[64]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[65]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[66]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[67]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[68]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[69]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[70]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[71]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[72]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[73]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[74]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[75]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[76]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[77]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[78]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[79]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[80]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[81]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[82]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[83]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[84]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[85]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_user_t[86]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[39]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[40]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[41]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[42]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[43]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[44]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[45]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[46]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[47]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[48]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[49]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[50]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[51]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[52]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[53]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[54]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[55]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[56]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[57]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[58]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[59]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[60]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[61]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[62]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[63]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[64]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[65]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[66]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[67]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[68]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[69]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[70]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[71]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[72]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[73]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[74]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[75]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[76]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[77]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[78]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[79]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[80]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[81]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[82]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[83]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[84]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[85]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
    //
    if (enToggle_past) begin
      cover(userBits_t[86]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 205:31]
    end
  end
endmodule
module PTERequestFilter(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input         io_out_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output        io_out_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input         io_out_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input  [63:0] io_out_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input         io_u // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
  wire  isLegal = |(io_in_req_bits_addr >= 32'h80000000); // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  _hasInflight_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [7:0] _io_in_resp_bits_rdata_T = {3'h7,io_u,4'hf}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 570:33]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  hasInflight_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
  wire  hasInflight_t = hasInflight ^ hasInflight_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
  wire  toggle_7419_clock;
  wire  toggle_7419_reset;
  wire  toggle_7419_valid;
  reg  toggle_7419_valid_reg;
  GEN_w1_toggle #(.COVER_INDEX(7419)) toggle_7419 (
    .clock(toggle_7419_clock),
    .reset(toggle_7419_reset),
    .valid(toggle_7419_valid)
  );
  assign io_in_req_ready = isLegal ? io_out_req_ready : ~hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 562:25]
  assign io_in_resp_valid = ~io_out_resp_valid & hasInflight | io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10 566:44 567:22]
  assign io_in_resp_bits_rdata = ~io_out_resp_valid & hasInflight ? {{56'd0}, _io_in_resp_bits_rdata_T} :
    io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10 566:44 570:27]
  assign io_out_req_valid = io_in_req_valid & isLegal; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 561:39]
  assign io_out_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10]
  assign io_out_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10]
  assign io_out_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10]
  assign toggle_7419_clock = clock;
  assign toggle_7419_reset = reset;
  assign toggle_7419_valid = hasInflight ^ toggle_7419_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
      hasInflight <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
    end else if (~io_out_resp_valid & hasInflight) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 566:44]
      hasInflight <= 1'h0;
    end else begin
      hasInflight <= _hasInflight_T & ~isLegal; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 564:15]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    hasInflight_p <= hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
    toggle_7419_valid_reg <= hasInflight;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  hasInflight = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  hasInflight_p = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  toggle_7419_valid_reg = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(hasInflight_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
    end
  end
endmodule
module Cache_fake(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [86:0] io_in_req_bits_user, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_in_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [86:0] io_in_resp_bits_user, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [1:0]  io_flush, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_out_mem_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_out_mem_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [31:0] io_out_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_out_mem_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_out_mem_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [63:0] io_out_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_mmio_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_mmio_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_mmio_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_mmio_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [63:0] io_mmio_resp_bits_rdata // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [95:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [95:0] _RAND_22;
  reg [95:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
  wire [31:0] _ismmio_T = io_in_req_bits_addr ^ 32'h30000000; // @[src/main/scala/nutcore/NutCore.scala 114:11]
  wire  _ismmio_T_2 = _ismmio_T[31:28] == 4'h0; // @[src/main/scala/nutcore/NutCore.scala 114:44]
  wire [31:0] _ismmio_T_3 = io_in_req_bits_addr ^ 32'h40000000; // @[src/main/scala/nutcore/NutCore.scala 114:11]
  wire  _ismmio_T_5 = _ismmio_T_3[31:30] == 2'h0; // @[src/main/scala/nutcore/NutCore.scala 114:44]
  wire  ismmio = _ismmio_T_2 | _ismmio_T_5; // @[src/main/scala/nutcore/NutCore.scala 115:15]
  wire  _ismmioRec_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  ismmioRec; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
  reg  needFlush; // @[src/main/scala/nutcore/mem/Cache.scala 566:26]
  wire  _GEN_1 = io_flush[0] & state != 3'h0 | needFlush; // @[src/main/scala/nutcore/mem/Cache.scala 566:26 567:{44,56}]
  wire  _alreadyOutFire_T = io_in_resp_ready & io_in_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
  wire  _GEN_3 = _alreadyOutFire_T | alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 570:{33,33,33}]
  wire  _T_11 = io_out_mem_req_ready & io_out_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_13 = io_out_mem_resp_ready & io_out_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _GEN_6 = _T_13 ? 3'h5 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 581:{37,45}]
  wire  _T_15 = io_mmio_req_ready & io_mmio_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _GEN_7 = _T_15 ? 3'h4 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 584:{33,41}]
  wire  _T_17 = io_mmio_resp_ready & io_mmio_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _GEN_8 = _T_17 | alreadyOutFire ? 3'h5 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 587:{52,60}]
  wire [2:0] _GEN_9 = _alreadyOutFire_T | needFlush | alreadyOutFire ? 3'h0 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 590:{63,71}]
  wire [2:0] _GEN_10 = 3'h5 == state ? _GEN_9 : state; // @[src/main/scala/nutcore/mem/Cache.scala 572:18 558:22]
  wire [2:0] _GEN_11 = 3'h4 == state ? _GEN_8 : _GEN_10; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  wire [2:0] _GEN_12 = 3'h3 == state ? _GEN_7 : _GEN_11; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  reg [31:0] reqaddr; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
  reg [63:0] mmiordata; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
  reg [63:0] memrdata; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
  reg [86:0] memuser; // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [2:0] state_p; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
  wire [2:0] state_t = state ^ state_p; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
  wire  toggle_7420_clock;
  wire  toggle_7420_reset;
  wire [2:0] toggle_7420_valid;
  reg [2:0] toggle_7420_valid_reg;
  reg  ismmioRec_p; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
  wire  ismmioRec_t = ismmioRec ^ ismmioRec_p; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
  wire  toggle_7423_clock;
  wire  toggle_7423_reset;
  wire  toggle_7423_valid;
  reg  toggle_7423_valid_reg;
  reg  needFlush_p; // @[src/main/scala/nutcore/mem/Cache.scala 566:26]
  wire  needFlush_t = needFlush ^ needFlush_p; // @[src/main/scala/nutcore/mem/Cache.scala 566:26]
  wire  toggle_7424_clock;
  wire  toggle_7424_reset;
  wire  toggle_7424_valid;
  reg  toggle_7424_valid_reg;
  reg  alreadyOutFire_p; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
  wire  alreadyOutFire_t = alreadyOutFire ^ alreadyOutFire_p; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
  wire  toggle_7425_clock;
  wire  toggle_7425_reset;
  wire  toggle_7425_valid;
  reg  toggle_7425_valid_reg;
  reg [31:0] reqaddr_p; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
  wire [31:0] reqaddr_t = reqaddr ^ reqaddr_p; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
  wire  toggle_7426_clock;
  wire  toggle_7426_reset;
  wire [31:0] toggle_7426_valid;
  reg [31:0] toggle_7426_valid_reg;
  reg [63:0] mmiordata_p; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
  wire [63:0] mmiordata_t = mmiordata ^ mmiordata_p; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
  wire  toggle_7458_clock;
  wire  toggle_7458_reset;
  wire [63:0] toggle_7458_valid;
  reg [63:0] toggle_7458_valid_reg;
  reg [63:0] memrdata_p; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
  wire [63:0] memrdata_t = memrdata ^ memrdata_p; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
  wire  toggle_7522_clock;
  wire  toggle_7522_reset;
  wire [63:0] toggle_7522_valid;
  reg [63:0] toggle_7522_valid_reg;
  reg [86:0] memuser_p; // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
  wire [86:0] memuser_t = memuser ^ memuser_p; // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
  wire  toggle_7586_clock;
  wire  toggle_7586_reset;
  wire [86:0] toggle_7586_valid;
  reg [86:0] toggle_7586_valid_reg;
  GEN_w3_toggle #(.COVER_INDEX(7420)) toggle_7420 (
    .clock(toggle_7420_clock),
    .reset(toggle_7420_reset),
    .valid(toggle_7420_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(7423)) toggle_7423 (
    .clock(toggle_7423_clock),
    .reset(toggle_7423_reset),
    .valid(toggle_7423_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(7424)) toggle_7424 (
    .clock(toggle_7424_clock),
    .reset(toggle_7424_reset),
    .valid(toggle_7424_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(7425)) toggle_7425 (
    .clock(toggle_7425_clock),
    .reset(toggle_7425_reset),
    .valid(toggle_7425_valid)
  );
  GEN_w32_toggle #(.COVER_INDEX(7426)) toggle_7426 (
    .clock(toggle_7426_clock),
    .reset(toggle_7426_reset),
    .valid(toggle_7426_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(7458)) toggle_7458 (
    .clock(toggle_7458_clock),
    .reset(toggle_7458_reset),
    .valid(toggle_7458_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(7522)) toggle_7522 (
    .clock(toggle_7522_clock),
    .reset(toggle_7522_reset),
    .valid(toggle_7522_valid)
  );
  GEN_w87_toggle #(.COVER_INDEX(7586)) toggle_7586 (
    .clock(toggle_7586_clock),
    .reset(toggle_7586_reset),
    .valid(toggle_7586_valid)
  );
  assign io_in_req_ready = state == 3'h0; // @[src/main/scala/nutcore/mem/Cache.scala 600:29]
  assign io_in_resp_valid = state == 3'h5 & ~needFlush; // @[src/main/scala/nutcore/mem/Cache.scala 601:47]
  assign io_in_resp_bits_rdata = ismmioRec ? mmiordata : memrdata; // @[src/main/scala/nutcore/mem/Cache.scala 608:31]
  assign io_in_resp_bits_user = memuser; // @[src/main/scala/nutcore/mem/Cache.scala 612:93]
  assign io_out_mem_req_valid = state == 3'h1; // @[src/main/scala/nutcore/mem/Cache.scala 617:34]
  assign io_out_mem_req_bits_addr = reqaddr; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_out_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 618:25]
  assign io_mmio_req_valid = state == 3'h3; // @[src/main/scala/nutcore/mem/Cache.scala 623:31]
  assign io_mmio_req_bits_addr = reqaddr; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_mmio_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 624:22]
  assign toggle_7420_clock = clock;
  assign toggle_7420_reset = reset;
  assign toggle_7420_valid = state ^ toggle_7420_valid_reg;
  assign toggle_7423_clock = clock;
  assign toggle_7423_reset = reset;
  assign toggle_7423_valid = ismmioRec ^ toggle_7423_valid_reg;
  assign toggle_7424_clock = clock;
  assign toggle_7424_reset = reset;
  assign toggle_7424_valid = needFlush ^ toggle_7424_valid_reg;
  assign toggle_7425_clock = clock;
  assign toggle_7425_reset = reset;
  assign toggle_7425_valid = alreadyOutFire ^ toggle_7425_valid_reg;
  assign toggle_7426_clock = clock;
  assign toggle_7426_reset = reset;
  assign toggle_7426_valid = reqaddr ^ toggle_7426_valid_reg;
  assign toggle_7458_clock = clock;
  assign toggle_7458_reset = reset;
  assign toggle_7458_valid = mmiordata ^ toggle_7458_valid_reg;
  assign toggle_7522_clock = clock;
  assign toggle_7522_reset = reset;
  assign toggle_7522_valid = memrdata ^ toggle_7522_valid_reg;
  assign toggle_7586_clock = clock;
  assign toggle_7586_reset = reset;
  assign toggle_7586_valid = memuser ^ toggle_7586_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
      state <= 3'h0; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      if (_ismmioRec_T & ~io_flush[0]) begin // @[src/main/scala/nutcore/mem/Cache.scala 575:47]
        if (ismmio) begin // @[src/main/scala/nutcore/mem/Cache.scala 575:61]
          state <= 3'h3;
        end else begin
          state <= 3'h1;
        end
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      if (_T_11) begin // @[src/main/scala/nutcore/mem/Cache.scala 578:36]
        state <= 3'h2; // @[src/main/scala/nutcore/mem/Cache.scala 578:44]
      end
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      state <= _GEN_6;
    end else begin
      state <= _GEN_12;
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
      ismmioRec <= ismmio; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 566:26]
      needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 566:26]
    end else if (state == 3'h0 & needFlush) begin // @[src/main/scala/nutcore/mem/Cache.scala 568:40]
      needFlush <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 568:52]
    end else begin
      needFlush <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 574:22]
    end else begin
      alreadyOutFire <= _GEN_3;
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
      reqaddr <= io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    if (_T_17) begin // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
      mmiordata <= io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    if (_T_13) begin // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
      memrdata <= io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
      memuser <= io_in_req_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    state_p <= state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
    toggle_7420_valid_reg <= state;
    ismmioRec_p <= ismmioRec; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
    toggle_7423_valid_reg <= ismmioRec;
    needFlush_p <= needFlush; // @[src/main/scala/nutcore/mem/Cache.scala 566:26]
    toggle_7424_valid_reg <= needFlush;
    alreadyOutFire_p <= alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
    toggle_7425_valid_reg <= alreadyOutFire;
    reqaddr_p <= reqaddr; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    toggle_7426_valid_reg <= reqaddr;
    mmiordata_p <= mmiordata; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    toggle_7458_valid_reg <= mmiordata;
    memrdata_p <= memrdata; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    toggle_7522_valid_reg <= memrdata;
    memuser_p <= memuser; // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    toggle_7586_valid_reg <= memuser;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  ismmioRec = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  needFlush = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  alreadyOutFire = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  reqaddr = _RAND_4[31:0];
  _RAND_5 = {2{`RANDOM}};
  mmiordata = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  memrdata = _RAND_6[63:0];
  _RAND_7 = {3{`RANDOM}};
  memuser = _RAND_7[86:0];
  _RAND_8 = {1{`RANDOM}};
  state_p = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  toggle_7420_valid_reg = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  ismmioRec_p = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  toggle_7423_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  needFlush_p = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  toggle_7424_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  alreadyOutFire_p = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  toggle_7425_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  reqaddr_p = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  toggle_7426_valid_reg = _RAND_17[31:0];
  _RAND_18 = {2{`RANDOM}};
  mmiordata_p = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  toggle_7458_valid_reg = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  memrdata_p = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  toggle_7522_valid_reg = _RAND_21[63:0];
  _RAND_22 = {3{`RANDOM}};
  memuser_p = _RAND_22[86:0];
  _RAND_23 = {3{`RANDOM}};
  toggle_7586_valid_reg = _RAND_23[86:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(state_t[0]); // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[1]); // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[2]); // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
    end
    //
    if (enToggle_past) begin
      cover(ismmioRec_t); // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
    end
    //
    if (enToggle_past) begin
      cover(needFlush_t); // @[src/main/scala/nutcore/mem/Cache.scala 566:26]
    end
    //
    if (enToggle_past) begin
      cover(alreadyOutFire_t); // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[0]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[1]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[2]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[3]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[4]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[5]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[6]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[7]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[8]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[9]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[10]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[11]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[12]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[13]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[14]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[15]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[16]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[17]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[18]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[19]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[20]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[21]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[22]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[23]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[24]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[25]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[26]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[27]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[28]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[29]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[30]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[31]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[0]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[1]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[2]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[3]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[4]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[5]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[6]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[7]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[8]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[9]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[10]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[11]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[12]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[13]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[14]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[15]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[16]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[17]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[18]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[19]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[20]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[21]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[22]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[23]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[24]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[25]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[26]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[27]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[28]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[29]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[30]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[31]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[32]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[33]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[34]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[35]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[36]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[37]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[38]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[39]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[40]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[41]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[42]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[43]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[44]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[45]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[46]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[47]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[48]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[49]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[50]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[51]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[52]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[53]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[54]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[55]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[56]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[57]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[58]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[59]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[60]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[61]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[62]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[63]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[0]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[1]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[2]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[3]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[4]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[5]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[6]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[7]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[8]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[9]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[10]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[11]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[12]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[13]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[14]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[15]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[16]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[17]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[18]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[19]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[20]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[21]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[22]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[23]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[24]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[25]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[26]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[27]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[28]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[29]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[30]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[31]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[32]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[33]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[34]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[35]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[36]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[37]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[38]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[39]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[40]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[41]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[42]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[43]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[44]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[45]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[46]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[47]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[48]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[49]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[50]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[51]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[52]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[53]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[54]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[55]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[56]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[57]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[58]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[59]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[60]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[61]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[62]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[63]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[0]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[1]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[2]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[3]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[4]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[5]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[6]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[7]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[8]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[9]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[10]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[11]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[12]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[13]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[14]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[15]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[16]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[17]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[18]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[19]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[20]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[21]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[22]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[23]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[24]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[25]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[26]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[27]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[28]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[29]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[30]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[31]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[32]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[33]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[34]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[35]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[36]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[37]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[38]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[39]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[40]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[41]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[42]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[43]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[44]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[45]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[46]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[47]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[48]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[49]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[50]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[51]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[52]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[53]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[54]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[55]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[56]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[57]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[58]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[59]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[60]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[61]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[62]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[63]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[64]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[65]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[66]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[67]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[68]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[69]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[70]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[71]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[72]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[73]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[74]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[75]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[76]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[77]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[78]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[79]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[80]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[81]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[82]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[83]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[84]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[85]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
    //
    if (enToggle_past) begin
      cover(memuser_t[86]); // @[src/main/scala/nutcore/mem/Cache.scala 611:26]
    end
  end
endmodule
module EmbeddedTLBExec_1(
  input          clock,
  input          reset,
  output         io_in_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_in_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [38:0]  io_in_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [2:0]   io_in_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [3:0]   io_in_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [7:0]   io_in_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [63:0]  io_in_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_out_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_out_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [31:0]  io_out_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [2:0]   io_out_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [3:0]   io_out_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [7:0]   io_out_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [63:0]  io_out_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_0, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_1, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_2, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [144:0] io_md_3, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_mdWrite_wen, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [3:0]   io_mdWrite_windex, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [3:0]   io_mdWrite_waymask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [144:0] io_mdWrite_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_mdReady, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_mem_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_mem_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [31:0]  io_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [3:0]   io_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output [63:0]  io_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_mem_resp_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_mem_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [63:0]  io_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [63:0]  io_satp, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input  [1:0]   io_pf_priviledgeMode, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_pf_status_sum, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          io_pf_status_mxr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_loadPF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_storePF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_laf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_pf_saf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  output         io_isFinish, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 221:14]
  input          lr_0,
  input          scInflight_0,
  input          ISAMO,
  input  [63:0]  lr_addr,
  output [55:0]  paddr_0,
  output         scIsSuccess_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] vpn_vpn0 = io_in_bits_addr[20:12]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:54]
  wire [8:0] vpn_vpn1 = io_in_bits_addr[29:21]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:54]
  wire [8:0] vpn_vpn2 = io_in_bits_addr[38:30]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 242:54]
  wire [43:0] satp_ppn = io_satp[43:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 244:30]
  wire [15:0] satp_asid = io_satp[59:44]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 244:30]
  wire [17:0] hitVec_hi = {vpn_vpn2,vpn_vpn1}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:201]
  wire [26:0] _hitVec_T_34 = {vpn_vpn2,vpn_vpn1,vpn_vpn0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:201]
  wire [26:0] _hitVec_T_35 = {9'h1ff,io_md_0[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_36 = _hitVec_T_35 & io_md_0[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_38 = _hitVec_T_35 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_39 = _hitVec_T_36 == _hitVec_T_38; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_40 = io_md_0[76] & io_md_0[117:102] == satp_asid & _hitVec_T_39; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [26:0] _hitVec_T_76 = {9'h1ff,io_md_1[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_77 = _hitVec_T_76 & io_md_1[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_79 = _hitVec_T_76 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_80 = _hitVec_T_77 == _hitVec_T_79; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_81 = io_md_1[76] & io_md_1[117:102] == satp_asid & _hitVec_T_80; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [26:0] _hitVec_T_117 = {9'h1ff,io_md_2[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_118 = _hitVec_T_117 & io_md_2[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_120 = _hitVec_T_117 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_121 = _hitVec_T_118 == _hitVec_T_120; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_122 = io_md_2[76] & io_md_2[117:102] == satp_asid & _hitVec_T_121; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [26:0] _hitVec_T_158 = {9'h1ff,io_md_3[101:84]}; // @[src/main/scala/nutcore/mem/TLB.scala 131:9]
  wire [26:0] _hitVec_T_159 = _hitVec_T_158 & io_md_3[144:118]; // @[src/main/scala/nutcore/mem/TLB.scala 131:37]
  wire [26:0] _hitVec_T_161 = _hitVec_T_158 & _hitVec_T_34; // @[src/main/scala/nutcore/mem/TLB.scala 131:84]
  wire  _hitVec_T_162 = _hitVec_T_159 == _hitVec_T_161; // @[src/main/scala/nutcore/mem/TLB.scala 131:48]
  wire  _hitVec_T_163 = io_md_3[76] & io_md_3[117:102] == satp_asid & _hitVec_T_162; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:132]
  wire [3:0] hitVec = {_hitVec_T_163,_hitVec_T_122,_hitVec_T_81,_hitVec_T_40}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 248:211]
  wire  _hit_T = |hitVec; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 249:35]
  wire  hit = io_in_valid & |hitVec; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 249:25]
  wire  miss = io_in_valid & ~_hit_T; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 250:26]
  reg [63:0] victimWaymask_lfsr; // @[src/main/scala/utils/LFSR64.scala 25:23]
  wire  victimWaymask_xor = victimWaymask_lfsr[0] ^ victimWaymask_lfsr[1] ^ victimWaymask_lfsr[3] ^ victimWaymask_lfsr[4
    ]; // @[src/main/scala/utils/LFSR64.scala 26:43]
  wire [63:0] _victimWaymask_lfsr_T_2 = {victimWaymask_xor,victimWaymask_lfsr[63:1]}; // @[src/main/scala/utils/LFSR64.scala 28:41]
  wire [3:0] victimWaymask = 4'h1 << victimWaymask_lfsr[1:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 252:42]
  wire [3:0] waymask = hit ? hitVec : victimWaymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:20]
  wire [144:0] _hitMeta_T_4 = waymask[0] ? io_md_0 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_5 = waymask[1] ? io_md_1 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_6 = waymask[2] ? io_md_2 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_7 = waymask[3] ? io_md_3 : 145'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_8 = _hitMeta_T_4 | _hitMeta_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_9 = _hitMeta_T_8 | _hitMeta_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [144:0] _hitMeta_T_10 = _hitMeta_T_9 | _hitMeta_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] hitMeta_flag = _hitMeta_T_10[83:76]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 262:70]
  wire [17:0] hitMeta_mask = _hitMeta_T_10[101:84]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 262:70]
  wire [43:0] hitData_ppn = _hitMeta_T_10[75:32]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 263:70]
  wire  hitFlag_r = hitMeta_flag[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_w = hitMeta_flag[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_x = hitMeta_flag[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_u = hitMeta_flag[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_a = hitMeta_flag[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire  hitFlag_d = hitMeta_flag[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 264:38]
  wire [7:0] _hitRefillFlag_T_1 = {io_in_bits_cmd[0],1'h1,6'h0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 269:26]
  wire  _hitCheck_T = io_pf_priviledgeMode == 2'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:62]
  wire  _hitCheck_T_5 = io_pf_priviledgeMode == 2'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:110]
  wire  _hitCheck_T_7 = ~io_pf_status_sum; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:137]
  wire  hitCheck = hit & ~(io_pf_priviledgeMode == 2'h0 & ~hitFlag_u) & ~(io_pf_priviledgeMode == 2'h1 & hitFlag_u & ~
    io_pf_status_sum); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 273:87]
  wire  hitADCheck = ~hitFlag_a | ~hitFlag_d & io_in_bits_cmd[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 274:31]
  wire  _hitExec_T_1 = hitCheck & ~hitADCheck; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 275:26]
  wire  hitLoad = _hitExec_T_1 & (hitFlag_r | io_pf_status_mxr & hitFlag_x); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 276:41]
  wire  hitStore = _hitExec_T_1 & hitFlag_w; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 277:42]
  reg  io_pf_loadPF_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:26]
  reg  io_pf_storePF_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 285:27]
  reg  io_pf_laf_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:23]
  reg  io_pf_saf_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:23]
  wire  _loadPF_T_5 = ~io_in_bits_cmd[0] & ~io_in_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _loadPF_T_7 = ~hitLoad & _loadPF_T_5 & hit; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:40]
  wire  _loadPF_T_8 = ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:50]
  reg [2:0] state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
  reg [1:0] level; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
  reg [63:0] memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
  reg [17:0] missMaskStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
  wire  memRdata_flag_v = io_mem_resp_bits_rdata[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_r = io_mem_resp_bits_rdata[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_w = io_mem_resp_bits_rdata[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_x = io_mem_resp_bits_rdata[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_u = io_mem_resp_bits_rdata[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_g = io_mem_resp_bits_rdata[5]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_a = io_mem_resp_bits_rdata[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire  memRdata_flag_d = io_mem_resp_bits_rdata[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire [43:0] memRdata_ppn = io_mem_resp_bits_rdata[53:10]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  wire [9:0] memRdata_reserved = io_mem_resp_bits_rdata[63:54]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
  reg [55:0] raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
  wire  _raddrCancel_T_3 = |(raddr >= 56'h80000000 & raddr < 56'h100000000); // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  raddrCancel = ~_raddrCancel_T_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 308:21]
  wire  _alreadyOutFire_T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  alreadyOutFire; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
  wire  _GEN_2 = _alreadyOutFire_T | alreadyOutFire; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:{33,33,33}]
  reg  missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
  wire [55:0] _raddr_T_1 = {satp_ppn,vpn_vpn2,3'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 89:8]
  wire  _T_10 = io_mem_req_ready & io_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _GEN_15 = raddrCancel ? 3'h5 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 343:32 344:59]
  wire  _GEN_16 = raddrCancel | missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 343:32 345:19 319:26]
  wire [7:0] _missflag_T = {memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,memRdata_flag_u,memRdata_flag_x,
    memRdata_flag_w,memRdata_flag_r,memRdata_flag_v}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_v = _missflag_T[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_r = _missflag_T[1]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_w = _missflag_T[2]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_x = _missflag_T[3]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_u = _missflag_T[4]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_g = _missflag_T[5]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_a = _missflag_T[6]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  missflag_d = _missflag_T[7]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 350:44]
  wire  _T_12 = io_mem_resp_ready & io_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_15 = level == 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:58]
  wire  _T_16 = level == 2'h2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:73]
  wire  _T_21 = ~missflag_r & missflag_w; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:44]
  wire  _loadPF_T_16 = _loadPF_T_5 & _loadPF_T_8; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 360:38]
  wire  _storePF_T_15 = io_in_bits_cmd[0] | ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 361:40]
  wire [8:0] _raddr_T_3 = _T_15 ? vpn_vpn1 : vpn_vpn0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 369:50]
  wire [55:0] _raddr_T_5 = {memRdata_ppn,_raddr_T_3,3'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 89:8]
  wire  is_reserved = memRdata_reserved != 10'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 370:49]
  wire [2:0] _GEN_22 = is_reserved ? 3'h5 : 3'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 368:19 371:32 377:23]
  wire  _GEN_23 = is_reserved ? _loadPF_T_16 : ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 371:32 378:24]
  wire  _GEN_24 = is_reserved ? _storePF_T_15 : ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 371:32 379:25]
  wire [2:0] _GEN_25 = ~missflag_v | ~missflag_r & missflag_w ? 3'h5 : _GEN_22; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:60 357:73]
  wire  _GEN_26 = ~missflag_v | ~missflag_r & missflag_w ? _loadPF_T_5 & _loadPF_T_8 : _GEN_23; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:60 360:22]
  wire  _GEN_27 = ~missflag_v | ~missflag_r & missflag_w ? io_in_bits_cmd[0] | ISAMO : _GEN_24; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 356:60 361:23]
  wire [55:0] _GEN_28 = ~missflag_v | ~missflag_r & missflag_w ? raddr : _raddr_T_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18 356:60 369:19]
  wire [17:0] pg_mask = _T_16 ? 18'h1ff : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 384:28]
  wire [43:0] _GEN_60 = {{26'd0}, pg_mask}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:54]
  wire [43:0] _misaligned_T_1 = memRdata_ppn & _GEN_60; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:54]
  wire  misaligned = level[1] & |_misaligned_T_1 | is_reserved; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 385:76]
  wire  permCheck = missflag_v & ~(_hitCheck_T & ~missflag_u) & ~(_hitCheck_T_5 & missflag_u & _hitCheck_T_7); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 386:87]
  wire  permAD = ~missflag_a | ~missflag_d & io_in_bits_cmd[0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 388:36]
  wire  _permExec_T_5 = permCheck & ~_T_21 & ~permAD & ~misaligned; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 389:60]
  wire  permLoad = _permExec_T_5 & (missflag_r | io_pf_status_mxr & missflag_x); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 390:75]
  wire  permStore = _permExec_T_5 & missflag_w; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 391:76]
  wire [63:0] updateData = {56'h0,io_in_bits_cmd[0],7'h40}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 392:31]
  wire [7:0] _missRefillFlag_T_2 = {missflag_d,missflag_a,missflag_g,missflag_u,missflag_x,missflag_w,missflag_r,
    missflag_v}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 393:79]
  wire [7:0] _missRefillFlag_T_3 = _hitRefillFlag_T_1 | _missRefillFlag_T_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 393:68]
  wire [63:0] _memRespStore_T = io_mem_resp_bits_rdata | updateData; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 394:50]
  wire [2:0] _GEN_29 = ~permLoad & _loadPF_T_5 | ~permStore & io_in_bits_cmd[0] ? 3'h5 : 3'h4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 403:80 404:21 408:21]
  wire  _GEN_30 = ~permLoad & _loadPF_T_5 | ~permStore & io_in_bits_cmd[0] ? _loadPF_T_16 : ~hitLoad & _loadPF_T_5 & hit
     & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 403:80 405:22]
  wire  _GEN_31 = ~permLoad & _loadPF_T_5 | ~permStore & io_in_bits_cmd[0] ? _storePF_T_15 : ~hitStore & io_in_bits_cmd[
    0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 403:80 406:23]
  wire  _GEN_32 = ~permLoad & _loadPF_T_5 | ~permStore & io_in_bits_cmd[0] ? 1'h0 : 1'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 403:80 409:30]
  wire [17:0] _missMask_T_2 = _T_16 ? 18'h3fe00 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 412:59]
  wire [17:0] _missMask_T_3 = _T_15 ? 18'h0 : _missMask_T_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 412:26]
  wire [7:0] _GEN_33 = level != 2'h0 ? _missRefillFlag_T_3 : 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 393:26 305:32]
  wire [63:0] _GEN_34 = level != 2'h0 ? _memRespStore_T : memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 394:24 301:25]
  wire [2:0] _GEN_35 = level != 2'h0 ? _GEN_29 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 383:36]
  wire  _GEN_36 = level != 2'h0 ? _GEN_30 : ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 383:36]
  wire  _GEN_37 = level != 2'h0 ? _GEN_31 : ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 383:36]
  wire  _GEN_38 = level != 2'h0 & _GEN_32; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 383:36]
  wire [17:0] _GEN_39 = level != 2'h0 ? _missMask_T_3 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 412:20 302:26]
  wire [17:0] _GEN_48 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 18'h3ffff : _GEN_39; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26 355:82]
  wire [17:0] _GEN_67 = _T_12 ? _GEN_48 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26 351:33]
  wire [17:0] _GEN_95 = 3'h2 == state ? _GEN_67 : 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 302:26]
  wire [17:0] _GEN_110 = 3'h1 == state ? 18'h3ffff : _GEN_95; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 302:26]
  wire [17:0] missMask = 3'h0 == state ? 18'h3ffff : _GEN_110; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 302:26]
  wire [17:0] _GEN_40 = level != 2'h0 ? missMask : missMaskStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 383:36 413:25 303:26]
  wire [2:0] _GEN_41 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_25 : _GEN_35; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:82]
  wire  _GEN_42 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_26 : _GEN_36; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:82]
  wire  _GEN_43 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_27 : _GEN_37; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 355:82]
  wire [55:0] _GEN_44 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? _GEN_28 : raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18 355:82]
  wire [7:0] _GEN_45 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 8'h0 : _GEN_33; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32 355:82]
  wire [63:0] _GEN_46 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? memRespStore : _GEN_34; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25 355:82]
  wire  _GEN_47 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? 1'h0 : _GEN_38; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 355:82]
  wire [17:0] _GEN_49 = ~(missflag_r | missflag_x) & (level == 2'h3 | level == 2'h2) ? missMaskStore : _GEN_40; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26 355:82]
  wire [1:0] _level_T_1 = level - 2'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 415:24]
  wire [2:0] _GEN_59 = _T_12 ? _GEN_41 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 351:33]
  wire  _GEN_61 = _T_12 ? _GEN_42 : ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 351:33]
  wire  _GEN_62 = _T_12 ? _GEN_43 : ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 351:33]
  wire  _GEN_66 = _T_12 & _GEN_47; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32 351:33]
  wire [1:0] _GEN_69 = _T_12 ? _level_T_1 : level; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33 415:15 299:22]
  wire [2:0] _GEN_70 = _T_10 ? 3'h4 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22 423:{38,46}]
  wire [2:0] _GEN_72 = io_isFinish | alreadyOutFire ? 3'h0 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 427:13 298:22]
  wire  _GEN_74 = io_isFinish | alreadyOutFire ? 1'h0 : missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 429:17 319:26]
  wire  _GEN_75 = io_isFinish | alreadyOutFire ? 1'h0 : _GEN_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 426:71 430:22]
  wire [2:0] _GEN_76 = 3'h5 == state ? 3'h0 : state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 434:13 298:22]
  wire  _GEN_77 = 3'h5 == state ? 1'h0 : missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 435:17 319:26]
  wire [2:0] _GEN_78 = 3'h4 == state ? _GEN_72 : _GEN_76; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_80 = 3'h4 == state ? _GEN_74 : _GEN_77; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_81 = 3'h4 == state ? _GEN_75 : _GEN_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire [2:0] _GEN_82 = 3'h3 == state ? _GEN_70 : _GEN_78; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_85 = 3'h3 == state ? missPTEAF : _GEN_80; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 319:26]
  wire  _GEN_86 = 3'h3 == state ? _GEN_2 : _GEN_81; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
  wire  _GEN_89 = 3'h2 == state ? _GEN_61 : ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 322:18]
  wire  _GEN_90 = 3'h2 == state ? _GEN_62 : ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 322:18]
  wire  _GEN_104 = 3'h1 == state ? ~hitLoad & _loadPF_T_5 & hit & ~ISAMO : _GEN_89; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 322:18]
  wire  _GEN_105 = 3'h1 == state ? ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO : _GEN_90; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 322:18]
  wire  _GEN_109 = 3'h1 == state ? 1'h0 : 3'h2 == state & _GEN_66; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 304:32]
  wire  loadPF = 3'h0 == state ? ~hitLoad & _loadPF_T_5 & hit & ~ISAMO : _GEN_104; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12 322:18]
  wire  storePF = 3'h0 == state ? ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO : _GEN_105; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13 322:18]
  wire  missMetaRefill = 3'h0 == state ? 1'h0 : _GEN_109; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18 304:32]
  wire  cmd = state == 3'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 440:23]
  wire  _T_45 = state == 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:82]
  reg  REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
  reg [3:0] REG_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:21]
  reg [3:0] REG_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:60]
  reg [26:0] REG_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
  reg [15:0] REG_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
  reg [17:0] REG_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
  reg [7:0] REG_6; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
  reg [43:0] REG_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
  reg [55:0] REG_8; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
  wire [168:0] _io_mdWrite_wdata_T = {REG_3,REG_4,REG_5,REG_6,REG_7,REG_8}; // @[src/main/scala/nutcore/mem/TLB.scala 220:22]
  wire [55:0] mdWriteAddr = {memRdata_ppn,12'h0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 451:24]
  wire  _mdMayHasAF_T_2 = mdWriteAddr >= 56'h40000000 & mdWriteAddr < 56'h40001000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_5 = mdWriteAddr >= 56'h80000000 & mdWriteAddr < 56'h100000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [1:0] _mdMayHasAF_T_6 = {_mdMayHasAF_T_5,_mdMayHasAF_T_2}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _mdMayHasAF_T_7 = |_mdMayHasAF_T_6; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  _mdMayHasAF_T_11 = mdWriteAddr >= 56'h38000000 & mdWriteAddr < 56'h38010000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_14 = mdWriteAddr >= 56'h3c000000 & mdWriteAddr < 56'h40000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_17 = mdWriteAddr >= 56'h40600000 & mdWriteAddr < 56'h40600010; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_20 = mdWriteAddr >= 56'h50000000 & mdWriteAddr < 56'h50400000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_23 = mdWriteAddr >= 56'h40001000 & mdWriteAddr < 56'h40001008; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _mdMayHasAF_T_29 = mdWriteAddr >= 56'h40002000 & mdWriteAddr < 56'h40003000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [7:0] _mdMayHasAF_T_33 = {_mdMayHasAF_T_5,_mdMayHasAF_T_29,_mdMayHasAF_T_2,_mdMayHasAF_T_23,_mdMayHasAF_T_20,
    _mdMayHasAF_T_17,_mdMayHasAF_T_14,_mdMayHasAF_T_11}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _mdMayHasAF_T_34 = |_mdMayHasAF_T_33; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  mdMayHasAF = ~_mdMayHasAF_T_7 | ~_mdMayHasAF_T_34 | ~_mdMayHasAF_T_34; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 452:84]
  reg  blockRefill; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
  wire [55:0] vaddr_ext = {24'h0,io_in_bits_addr[31:0]}; // @[src/main/scala/utils/BitUtils.scala 49:41]
  wire [55:0] _paddr_T = {hitData_ppn,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:24]
  wire [55:0] _paddr_T_2 = {26'h3ffffff,hitMeta_mask,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:49]
  wire [55:0] _paddr_T_3 = _paddr_T & _paddr_T_2; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [55:0] _paddr_T_4 = ~_paddr_T_2; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [55:0] _paddr_T_5 = vaddr_ext & _paddr_T_4; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [55:0] _paddr_T_6 = _paddr_T_3 | _paddr_T_5; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [55:0] _paddr_T_18 = {memRespStore[53:10],12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:24]
  wire [55:0] _paddr_T_20 = {26'h3ffffff,missMaskStore,12'h0}; // @[src/main/scala/nutcore/mem/TLB.scala 127:49]
  wire [55:0] _paddr_T_21 = _paddr_T_18 & _paddr_T_20; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [55:0] _paddr_T_22 = ~_paddr_T_20; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [55:0] _paddr_T_23 = vaddr_ext & _paddr_T_22; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [55:0] _paddr_T_24 = _paddr_T_21 | _paddr_T_23; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire  _T_59 = ~scInflight_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 476:12]
  wire [55:0] paddr = hit ? _paddr_T_6 : _paddr_T_24; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 461:15]
  wire [63:0] _GEN_71 = {{8'd0}, paddr}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 477:49]
  wire  _scIsSuccess_T_7 = hit | state == 3'h4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 477:81]
  wire  out_req_valid = io_in_valid & _scIsSuccess_T_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 484:35]
  wire  _ldReqAF_T_2 = paddr >= 56'h38000000 & paddr < 56'h38010000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_5 = paddr >= 56'h3c000000 & paddr < 56'h40000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_8 = paddr >= 56'h40600000 & paddr < 56'h40600010; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_11 = paddr >= 56'h50000000 & paddr < 56'h50400000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_14 = paddr >= 56'h40001000 & paddr < 56'h40001008; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_17 = paddr >= 56'h40000000 & paddr < 56'h40001000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_20 = paddr >= 56'h40002000 & paddr < 56'h40003000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire  _ldReqAF_T_23 = paddr >= 56'h80000000 & paddr < 56'h100000000; // @[src/main/scala/nutcore/NutCore.scala 70:41]
  wire [7:0] _ldReqAF_T_24 = {_ldReqAF_T_23,_ldReqAF_T_20,_ldReqAF_T_17,_ldReqAF_T_14,_ldReqAF_T_11,_ldReqAF_T_8,
    _ldReqAF_T_5,_ldReqAF_T_2}; // @[src/main/scala/nutcore/NutCore.scala 70:60]
  wire  _ldReqAF_T_25 = |_ldReqAF_T_24; // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  ldReqAF = out_req_valid & ~_ldReqAF_T_25; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 489:34]
  wire  loadAF = (ldReqAF | missPTEAF) & _loadPF_T_5 & _loadPF_T_8; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 491:54]
  wire  storeAF = ldReqAF & io_in_bits_cmd[0] | ldReqAF & _loadPF_T_5 & ISAMO | missPTEAF & _storePF_T_15; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 492:79]
  wire  _hasException_T = io_pf_loadPF | io_pf_storePF; // @[src/main/scala/nutcore/Bundle.scala 134:23]
  wire  _hasException_T_1 = io_pf_laf | io_pf_saf; // @[src/main/scala/nutcore/Bundle.scala 135:24]
  wire  _hasException_T_2 = _hasException_T | _hasException_T_1; // @[src/main/scala/nutcore/Bundle.scala 136:35]
  wire  hasException = _hasException_T_2 | loadPF | storePF | loadAF | storeAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 494:72]
  wire  _io_out_valid_T_5 = ~hasException; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 496:78]
  wire  scIsSuccess = _T_59 | lr_0 & lr_addr == _GEN_71 | ~(hit | state == 3'h4); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 477:60]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [63:0] victimWaymask_lfsr_p; // @[src/main/scala/utils/LFSR64.scala 25:23]
  wire [63:0] victimWaymask_lfsr_t = victimWaymask_lfsr ^ victimWaymask_lfsr_p; // @[src/main/scala/utils/LFSR64.scala 25:23]
  wire  toggle_7673_clock;
  wire  toggle_7673_reset;
  wire [63:0] toggle_7673_valid;
  reg [63:0] toggle_7673_valid_reg;
  reg  io_pf_loadPF_REG_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:26]
  wire  io_pf_loadPF_REG_t = io_pf_loadPF_REG ^ io_pf_loadPF_REG_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:26]
  wire  toggle_7737_clock;
  wire  toggle_7737_reset;
  wire  toggle_7737_valid;
  reg  toggle_7737_valid_reg;
  reg  io_pf_storePF_REG_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 285:27]
  wire  io_pf_storePF_REG_t = io_pf_storePF_REG ^ io_pf_storePF_REG_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 285:27]
  wire  toggle_7738_clock;
  wire  toggle_7738_reset;
  wire  toggle_7738_valid;
  reg  toggle_7738_valid_reg;
  reg  io_pf_laf_REG_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:23]
  wire  io_pf_laf_REG_t = io_pf_laf_REG ^ io_pf_laf_REG_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:23]
  wire  toggle_7739_clock;
  wire  toggle_7739_reset;
  wire  toggle_7739_valid;
  reg  toggle_7739_valid_reg;
  reg  io_pf_saf_REG_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:23]
  wire  io_pf_saf_REG_t = io_pf_saf_REG ^ io_pf_saf_REG_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:23]
  wire  toggle_7740_clock;
  wire  toggle_7740_reset;
  wire  toggle_7740_valid;
  reg  toggle_7740_valid_reg;
  reg [2:0] state_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
  wire [2:0] state_t = state ^ state_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
  wire  toggle_7741_clock;
  wire  toggle_7741_reset;
  wire [2:0] toggle_7741_valid;
  reg [2:0] toggle_7741_valid_reg;
  reg [1:0] level_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
  wire [1:0] level_t = level ^ level_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
  wire  toggle_7744_clock;
  wire  toggle_7744_reset;
  wire [1:0] toggle_7744_valid;
  reg [1:0] toggle_7744_valid_reg;
  reg [63:0] memRespStore_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
  wire [63:0] memRespStore_t = memRespStore ^ memRespStore_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
  wire  toggle_7746_clock;
  wire  toggle_7746_reset;
  wire [63:0] toggle_7746_valid;
  reg [63:0] toggle_7746_valid_reg;
  reg [17:0] missMaskStore_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
  wire [17:0] missMaskStore_t = missMaskStore ^ missMaskStore_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
  wire  toggle_7810_clock;
  wire  toggle_7810_reset;
  wire [17:0] toggle_7810_valid;
  reg [17:0] toggle_7810_valid_reg;
  reg [55:0] raddr_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
  wire [55:0] raddr_t = raddr ^ raddr_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
  wire  toggle_7828_clock;
  wire  toggle_7828_reset;
  wire [55:0] toggle_7828_valid;
  reg [55:0] toggle_7828_valid_reg;
  reg  alreadyOutFire_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
  wire  alreadyOutFire_t = alreadyOutFire ^ alreadyOutFire_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
  wire  toggle_7884_clock;
  wire  toggle_7884_reset;
  wire  toggle_7884_valid;
  reg  toggle_7884_valid_reg;
  reg  missPTEAF_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
  wire  missPTEAF_t = missPTEAF ^ missPTEAF_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
  wire  toggle_7885_clock;
  wire  toggle_7885_reset;
  wire  toggle_7885_valid;
  reg  toggle_7885_valid_reg;
  reg  REG_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
  wire  REG_t = REG ^ REG_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
  wire  toggle_7886_clock;
  wire  toggle_7886_reset;
  wire  toggle_7886_valid;
  reg  toggle_7886_valid_reg;
  reg [3:0] REG_1_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:21]
  wire [3:0] REG_1_t = REG_1 ^ REG_1_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:21]
  wire  toggle_7887_clock;
  wire  toggle_7887_reset;
  wire [3:0] toggle_7887_valid;
  reg [3:0] toggle_7887_valid_reg;
  reg [3:0] REG_2_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:60]
  wire [3:0] REG_2_t = REG_2 ^ REG_2_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:60]
  wire  toggle_7891_clock;
  wire  toggle_7891_reset;
  wire [3:0] toggle_7891_valid;
  reg [3:0] toggle_7891_valid_reg;
  reg [26:0] REG_3_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
  wire [26:0] REG_3_t = REG_3 ^ REG_3_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
  wire  toggle_7895_clock;
  wire  toggle_7895_reset;
  wire [26:0] toggle_7895_valid;
  reg [26:0] toggle_7895_valid_reg;
  reg [15:0] REG_4_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
  wire [15:0] REG_4_t = REG_4 ^ REG_4_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
  wire  toggle_7922_clock;
  wire  toggle_7922_reset;
  wire [15:0] toggle_7922_valid;
  reg [15:0] toggle_7922_valid_reg;
  reg [17:0] REG_5_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
  wire [17:0] REG_5_t = REG_5 ^ REG_5_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
  wire  toggle_7938_clock;
  wire  toggle_7938_reset;
  wire [17:0] toggle_7938_valid;
  reg [17:0] toggle_7938_valid_reg;
  reg [7:0] REG_6_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
  wire [7:0] REG_6_t = REG_6 ^ REG_6_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
  wire  toggle_7956_clock;
  wire  toggle_7956_reset;
  wire [7:0] toggle_7956_valid;
  reg [7:0] toggle_7956_valid_reg;
  reg [43:0] REG_7_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
  wire [43:0] REG_7_t = REG_7 ^ REG_7_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
  wire  toggle_7964_clock;
  wire  toggle_7964_reset;
  wire [43:0] toggle_7964_valid;
  reg [43:0] toggle_7964_valid_reg;
  reg [55:0] REG_8_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
  wire [55:0] REG_8_t = REG_8 ^ REG_8_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
  wire  toggle_8008_clock;
  wire  toggle_8008_reset;
  wire [55:0] toggle_8008_valid;
  reg [55:0] toggle_8008_valid_reg;
  reg  blockRefill_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
  wire  blockRefill_t = blockRefill ^ blockRefill_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
  wire  toggle_8064_clock;
  wire  toggle_8064_reset;
  wire  toggle_8064_valid;
  reg  toggle_8064_valid_reg;
  GEN_w64_toggle #(.COVER_INDEX(7673)) toggle_7673 (
    .clock(toggle_7673_clock),
    .reset(toggle_7673_reset),
    .valid(toggle_7673_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(7737)) toggle_7737 (
    .clock(toggle_7737_clock),
    .reset(toggle_7737_reset),
    .valid(toggle_7737_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(7738)) toggle_7738 (
    .clock(toggle_7738_clock),
    .reset(toggle_7738_reset),
    .valid(toggle_7738_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(7739)) toggle_7739 (
    .clock(toggle_7739_clock),
    .reset(toggle_7739_reset),
    .valid(toggle_7739_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(7740)) toggle_7740 (
    .clock(toggle_7740_clock),
    .reset(toggle_7740_reset),
    .valid(toggle_7740_valid)
  );
  GEN_w3_toggle #(.COVER_INDEX(7741)) toggle_7741 (
    .clock(toggle_7741_clock),
    .reset(toggle_7741_reset),
    .valid(toggle_7741_valid)
  );
  GEN_w2_toggle #(.COVER_INDEX(7744)) toggle_7744 (
    .clock(toggle_7744_clock),
    .reset(toggle_7744_reset),
    .valid(toggle_7744_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(7746)) toggle_7746 (
    .clock(toggle_7746_clock),
    .reset(toggle_7746_reset),
    .valid(toggle_7746_valid)
  );
  GEN_w18_toggle #(.COVER_INDEX(7810)) toggle_7810 (
    .clock(toggle_7810_clock),
    .reset(toggle_7810_reset),
    .valid(toggle_7810_valid)
  );
  GEN_w56_toggle #(.COVER_INDEX(7828)) toggle_7828 (
    .clock(toggle_7828_clock),
    .reset(toggle_7828_reset),
    .valid(toggle_7828_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(7884)) toggle_7884 (
    .clock(toggle_7884_clock),
    .reset(toggle_7884_reset),
    .valid(toggle_7884_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(7885)) toggle_7885 (
    .clock(toggle_7885_clock),
    .reset(toggle_7885_reset),
    .valid(toggle_7885_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(7886)) toggle_7886 (
    .clock(toggle_7886_clock),
    .reset(toggle_7886_reset),
    .valid(toggle_7886_valid)
  );
  GEN_w4_toggle #(.COVER_INDEX(7887)) toggle_7887 (
    .clock(toggle_7887_clock),
    .reset(toggle_7887_reset),
    .valid(toggle_7887_valid)
  );
  GEN_w4_toggle #(.COVER_INDEX(7891)) toggle_7891 (
    .clock(toggle_7891_clock),
    .reset(toggle_7891_reset),
    .valid(toggle_7891_valid)
  );
  GEN_w27_toggle #(.COVER_INDEX(7895)) toggle_7895 (
    .clock(toggle_7895_clock),
    .reset(toggle_7895_reset),
    .valid(toggle_7895_valid)
  );
  GEN_w16_toggle #(.COVER_INDEX(7922)) toggle_7922 (
    .clock(toggle_7922_clock),
    .reset(toggle_7922_reset),
    .valid(toggle_7922_valid)
  );
  GEN_w18_toggle #(.COVER_INDEX(7938)) toggle_7938 (
    .clock(toggle_7938_clock),
    .reset(toggle_7938_reset),
    .valid(toggle_7938_valid)
  );
  GEN_w8_toggle #(.COVER_INDEX(7956)) toggle_7956 (
    .clock(toggle_7956_clock),
    .reset(toggle_7956_reset),
    .valid(toggle_7956_valid)
  );
  GEN_w44_toggle #(.COVER_INDEX(7964)) toggle_7964 (
    .clock(toggle_7964_clock),
    .reset(toggle_7964_reset),
    .valid(toggle_7964_valid)
  );
  GEN_w56_toggle #(.COVER_INDEX(8008)) toggle_8008 (
    .clock(toggle_8008_clock),
    .reset(toggle_8008_reset),
    .valid(toggle_8008_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(8064)) toggle_8064 (
    .clock(toggle_8064_clock),
    .reset(toggle_8064_reset),
    .valid(toggle_8064_valid)
  );
  assign io_in_ready = io_out_ready & _T_45 & ~miss & io_mdReady & _io_out_valid_T_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 498:86]
  assign io_out_valid = out_req_valid & ~hasException & scIsSuccess; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 496:92]
  assign io_out_bits_addr = paddr[31:0]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 483:20]
  assign io_out_bits_size = io_in_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 482:15]
  assign io_out_bits_cmd = io_in_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 482:15]
  assign io_out_bits_wmask = io_in_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 482:15]
  assign io_out_bits_wdata = io_in_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 482:15]
  assign io_mdWrite_wen = blockRefill ? 1'h0 : REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 454:22 455:20 src/main/scala/nutcore/mem/TLB.scala 217:14]
  assign io_mdWrite_windex = REG_1; // @[src/main/scala/nutcore/mem/TLB.scala 218:17]
  assign io_mdWrite_waymask = REG_2; // @[src/main/scala/nutcore/mem/TLB.scala 219:18]
  assign io_mdWrite_wdata = _io_mdWrite_wdata_T[144:0]; // @[src/main/scala/nutcore/mem/TLB.scala 220:16]
  assign io_mem_req_valid = (state == 3'h1 | cmd) & ~raddrCancel; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 442:85]
  assign io_mem_req_bits_addr = raddr[31:0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_mem_req_bits_cmd = {{3'd0}, cmd}; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 441:138]
  assign io_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 443:21]
  assign io_pf_loadPF = io_pf_loadPF_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:16]
  assign io_pf_storePF = io_pf_storePF_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 285:17]
  assign io_pf_laf = io_pf_laf_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:13]
  assign io_pf_saf = io_pf_saf_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:13]
  assign io_isFinish = _alreadyOutFire_T | _hasException_T_2 | ~scIsSuccess; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 502:54]
  assign paddr_0 = paddr;
  assign scIsSuccess_0 = scIsSuccess;
  assign toggle_7673_clock = clock;
  assign toggle_7673_reset = reset;
  assign toggle_7673_valid = victimWaymask_lfsr ^ toggle_7673_valid_reg;
  assign toggle_7737_clock = clock;
  assign toggle_7737_reset = reset;
  assign toggle_7737_valid = io_pf_loadPF_REG ^ toggle_7737_valid_reg;
  assign toggle_7738_clock = clock;
  assign toggle_7738_reset = reset;
  assign toggle_7738_valid = io_pf_storePF_REG ^ toggle_7738_valid_reg;
  assign toggle_7739_clock = clock;
  assign toggle_7739_reset = reset;
  assign toggle_7739_valid = io_pf_laf_REG ^ toggle_7739_valid_reg;
  assign toggle_7740_clock = clock;
  assign toggle_7740_reset = reset;
  assign toggle_7740_valid = io_pf_saf_REG ^ toggle_7740_valid_reg;
  assign toggle_7741_clock = clock;
  assign toggle_7741_reset = reset;
  assign toggle_7741_valid = state ^ toggle_7741_valid_reg;
  assign toggle_7744_clock = clock;
  assign toggle_7744_reset = reset;
  assign toggle_7744_valid = level ^ toggle_7744_valid_reg;
  assign toggle_7746_clock = clock;
  assign toggle_7746_reset = reset;
  assign toggle_7746_valid = memRespStore ^ toggle_7746_valid_reg;
  assign toggle_7810_clock = clock;
  assign toggle_7810_reset = reset;
  assign toggle_7810_valid = missMaskStore ^ toggle_7810_valid_reg;
  assign toggle_7828_clock = clock;
  assign toggle_7828_reset = reset;
  assign toggle_7828_valid = raddr ^ toggle_7828_valid_reg;
  assign toggle_7884_clock = clock;
  assign toggle_7884_reset = reset;
  assign toggle_7884_valid = alreadyOutFire ^ toggle_7884_valid_reg;
  assign toggle_7885_clock = clock;
  assign toggle_7885_reset = reset;
  assign toggle_7885_valid = missPTEAF ^ toggle_7885_valid_reg;
  assign toggle_7886_clock = clock;
  assign toggle_7886_reset = reset;
  assign toggle_7886_valid = REG ^ toggle_7886_valid_reg;
  assign toggle_7887_clock = clock;
  assign toggle_7887_reset = reset;
  assign toggle_7887_valid = REG_1 ^ toggle_7887_valid_reg;
  assign toggle_7891_clock = clock;
  assign toggle_7891_reset = reset;
  assign toggle_7891_valid = REG_2 ^ toggle_7891_valid_reg;
  assign toggle_7895_clock = clock;
  assign toggle_7895_reset = reset;
  assign toggle_7895_valid = REG_3 ^ toggle_7895_valid_reg;
  assign toggle_7922_clock = clock;
  assign toggle_7922_reset = reset;
  assign toggle_7922_valid = REG_4 ^ toggle_7922_valid_reg;
  assign toggle_7938_clock = clock;
  assign toggle_7938_reset = reset;
  assign toggle_7938_valid = REG_5 ^ toggle_7938_valid_reg;
  assign toggle_7956_clock = clock;
  assign toggle_7956_reset = reset;
  assign toggle_7956_valid = REG_6 ^ toggle_7956_valid_reg;
  assign toggle_7964_clock = clock;
  assign toggle_7964_reset = reset;
  assign toggle_7964_valid = REG_7 ^ toggle_7964_valid_reg;
  assign toggle_8008_clock = clock;
  assign toggle_8008_reset = reset;
  assign toggle_8008_valid = REG_8 ^ toggle_8008_valid_reg;
  assign toggle_8064_clock = clock;
  assign toggle_8064_reset = reset;
  assign toggle_8064_valid = blockRefill ^ toggle_8064_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/LFSR64.scala 25:23]
      victimWaymask_lfsr <= 64'h1234567887654321; // @[src/main/scala/utils/LFSR64.scala 25:23]
    end else if (victimWaymask_lfsr == 64'h0) begin // @[src/main/scala/utils/LFSR64.scala 28:18]
      victimWaymask_lfsr <= 64'h1;
    end else begin
      victimWaymask_lfsr <= _victimWaymask_lfsr_T_2;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:26]
      io_pf_loadPF_REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:26]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      io_pf_loadPF_REG <= ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      io_pf_loadPF_REG <= ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      io_pf_loadPF_REG <= _GEN_61;
    end else begin
      io_pf_loadPF_REG <= ~hitLoad & _loadPF_T_5 & hit & ~ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 292:12]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 285:27]
      io_pf_storePF_REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 285:27]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      io_pf_storePF_REG <= ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      io_pf_storePF_REG <= ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      io_pf_storePF_REG <= _GEN_62;
    end else begin
      io_pf_storePF_REG <= ~hitStore & io_in_bits_cmd[0] & hit | _loadPF_T_7 & ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 293:13]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:23]
      io_pf_laf_REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:23]
    end else begin
      io_pf_laf_REG <= loadAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:23]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:23]
      io_pf_saf_REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:23]
    end else begin
      io_pf_saf_REG <= storeAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:23]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
      state <= 3'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        state <= 3'h1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 329:15]
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (_T_10) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 341:38]
        state <= 3'h2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 342:15]
      end else begin
        state <= _GEN_15;
      end
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      state <= _GEN_59;
    end else begin
      state <= _GEN_82;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
      level <= 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        level <= 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 331:15]
      end
    end else if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        level <= _GEN_69;
      end
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
          if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
            memRespStore <= _GEN_46;
          end
        end
      end
    end
    if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
          if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
            missMaskStore <= _GEN_49;
          end
        end
      end
    end
    if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        raddr <= _raddr_T_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 330:15]
      end
    end else if (!(3'h1 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
          raddr <= _GEN_44;
        end
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (miss) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 328:37]
        alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 333:24]
      end else begin
        alreadyOutFire <= _GEN_2;
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      alreadyOutFire <= _GEN_2;
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      alreadyOutFire <= _GEN_2;
    end else begin
      alreadyOutFire <= _GEN_86;
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
      missPTEAF <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
    end else if (!(3'h0 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        if (!(_T_10)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 341:38]
          missPTEAF <= _GEN_16;
        end
      end else if (!(3'h2 == state)) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
        missPTEAF <= _GEN_85;
      end
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
      REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 304:32]
    end else begin
      REG <= 3'h2 == state & _GEN_66;
    end
    REG_1 <= io_in_bits_addr[15:12]; // @[src/main/scala/nutcore/mem/TLB.scala 203:19]
    if (hit) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 253:20]
      REG_2 <= hitVec;
    end else begin
      REG_2 <= victimWaymask;
    end
    REG_3 <= {hitVec_hi,vpn_vpn0}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:89]
    REG_4 <= io_satp[59:44]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 244:30]
    if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
        REG_5 <= _GEN_48;
      end else begin
        REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
      end
    end else begin
      REG_5 <= 18'h3ffff; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 302:26]
    end
    if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 322:18]
      if (_T_12) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 351:33]
        REG_6 <= _GEN_45;
      end else begin
        REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
      end
    end else begin
      REG_6 <= 8'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 305:32]
    end
    REG_7 <= io_mem_resp_bits_rdata[53:10]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 306:49]
    REG_8 <= raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:27]
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
      blockRefill <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
    end else begin
      blockRefill <= missMetaRefill & mdMayHasAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~scInflight_0 | ~io_in_valid | io_in_bits_cmd[0])) begin
          $fwrite(32'h80000002,
            "Assertion failed: SC is inflight but TLB receives a read request\n    at EmbeddedTLB.scala:476 assert(!scInflight || !io.in.valid || req.isWrite(), \"SC is inflight but TLB receives a read request\")\n"
            ); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 476:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    victimWaymask_lfsr_p <= victimWaymask_lfsr; // @[src/main/scala/utils/LFSR64.scala 25:23]
    toggle_7673_valid_reg <= victimWaymask_lfsr;
    io_pf_loadPF_REG_p <= io_pf_loadPF_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:26]
    toggle_7737_valid_reg <= io_pf_loadPF_REG;
    io_pf_storePF_REG_p <= io_pf_storePF_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 285:27]
    toggle_7738_valid_reg <= io_pf_storePF_REG;
    io_pf_laf_REG_p <= io_pf_laf_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:23]
    toggle_7739_valid_reg <= io_pf_laf_REG;
    io_pf_saf_REG_p <= io_pf_saf_REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:23]
    toggle_7740_valid_reg <= io_pf_saf_REG;
    state_p <= state; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
    toggle_7741_valid_reg <= state;
    level_p <= level; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
    toggle_7744_valid_reg <= level;
    memRespStore_p <= memRespStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    toggle_7746_valid_reg <= memRespStore;
    missMaskStore_p <= missMaskStore; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    toggle_7810_valid_reg <= missMaskStore;
    raddr_p <= raddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    toggle_7828_valid_reg <= raddr;
    alreadyOutFire_p <= alreadyOutFire; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
    toggle_7884_valid_reg <= alreadyOutFire;
    missPTEAF_p <= missPTEAF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
    toggle_7885_valid_reg <= missPTEAF;
    REG_p <= REG; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
    toggle_7886_valid_reg <= REG;
    REG_1_p <= REG_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:21]
    toggle_7887_valid_reg <= REG_1;
    REG_2_p <= REG_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:60]
    toggle_7891_valid_reg <= REG_2;
    REG_3_p <= REG_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    toggle_7895_valid_reg <= REG_3;
    REG_4_p <= REG_4; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    toggle_7922_valid_reg <= REG_4;
    REG_5_p <= REG_5; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    toggle_7938_valid_reg <= REG_5;
    REG_6_p <= REG_6; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
    toggle_7956_valid_reg <= REG_6;
    REG_7_p <= REG_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    toggle_7964_valid_reg <= REG_7;
    REG_8_p <= REG_8; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    toggle_8008_valid_reg <= REG_8;
    blockRefill_p <= blockRefill; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
    toggle_8064_valid_reg <= blockRefill;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  victimWaymask_lfsr = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  io_pf_loadPF_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_pf_storePF_REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  io_pf_laf_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_pf_saf_REG = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  level = _RAND_6[1:0];
  _RAND_7 = {2{`RANDOM}};
  memRespStore = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  missMaskStore = _RAND_8[17:0];
  _RAND_9 = {2{`RANDOM}};
  raddr = _RAND_9[55:0];
  _RAND_10 = {1{`RANDOM}};
  alreadyOutFire = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  missPTEAF = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  REG = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  REG_1 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  REG_2 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  REG_3 = _RAND_15[26:0];
  _RAND_16 = {1{`RANDOM}};
  REG_4 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  REG_5 = _RAND_17[17:0];
  _RAND_18 = {1{`RANDOM}};
  REG_6 = _RAND_18[7:0];
  _RAND_19 = {2{`RANDOM}};
  REG_7 = _RAND_19[43:0];
  _RAND_20 = {2{`RANDOM}};
  REG_8 = _RAND_20[55:0];
  _RAND_21 = {1{`RANDOM}};
  blockRefill = _RAND_21[0:0];
  _RAND_22 = {2{`RANDOM}};
  victimWaymask_lfsr_p = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  toggle_7673_valid_reg = _RAND_23[63:0];
  _RAND_24 = {1{`RANDOM}};
  io_pf_loadPF_REG_p = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  toggle_7737_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  io_pf_storePF_REG_p = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  toggle_7738_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  io_pf_laf_REG_p = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  toggle_7739_valid_reg = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  io_pf_saf_REG_p = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  toggle_7740_valid_reg = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  state_p = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  toggle_7741_valid_reg = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  level_p = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  toggle_7744_valid_reg = _RAND_35[1:0];
  _RAND_36 = {2{`RANDOM}};
  memRespStore_p = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  toggle_7746_valid_reg = _RAND_37[63:0];
  _RAND_38 = {1{`RANDOM}};
  missMaskStore_p = _RAND_38[17:0];
  _RAND_39 = {1{`RANDOM}};
  toggle_7810_valid_reg = _RAND_39[17:0];
  _RAND_40 = {2{`RANDOM}};
  raddr_p = _RAND_40[55:0];
  _RAND_41 = {2{`RANDOM}};
  toggle_7828_valid_reg = _RAND_41[55:0];
  _RAND_42 = {1{`RANDOM}};
  alreadyOutFire_p = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  toggle_7884_valid_reg = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  missPTEAF_p = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  toggle_7885_valid_reg = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  REG_p = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  toggle_7886_valid_reg = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  REG_1_p = _RAND_48[3:0];
  _RAND_49 = {1{`RANDOM}};
  toggle_7887_valid_reg = _RAND_49[3:0];
  _RAND_50 = {1{`RANDOM}};
  REG_2_p = _RAND_50[3:0];
  _RAND_51 = {1{`RANDOM}};
  toggle_7891_valid_reg = _RAND_51[3:0];
  _RAND_52 = {1{`RANDOM}};
  REG_3_p = _RAND_52[26:0];
  _RAND_53 = {1{`RANDOM}};
  toggle_7895_valid_reg = _RAND_53[26:0];
  _RAND_54 = {1{`RANDOM}};
  REG_4_p = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  toggle_7922_valid_reg = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  REG_5_p = _RAND_56[17:0];
  _RAND_57 = {1{`RANDOM}};
  toggle_7938_valid_reg = _RAND_57[17:0];
  _RAND_58 = {1{`RANDOM}};
  REG_6_p = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  toggle_7956_valid_reg = _RAND_59[7:0];
  _RAND_60 = {2{`RANDOM}};
  REG_7_p = _RAND_60[43:0];
  _RAND_61 = {2{`RANDOM}};
  toggle_7964_valid_reg = _RAND_61[43:0];
  _RAND_62 = {2{`RANDOM}};
  REG_8_p = _RAND_62[55:0];
  _RAND_63 = {2{`RANDOM}};
  toggle_8008_valid_reg = _RAND_63[55:0];
  _RAND_64 = {1{`RANDOM}};
  blockRefill_p = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  toggle_8064_valid_reg = _RAND_65[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~scInflight_0 | ~io_in_valid | io_in_bits_cmd[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 476:11]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[0]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[1]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[2]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[3]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[4]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[5]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[6]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[7]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[8]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[9]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[10]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[11]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[12]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[13]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[14]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[15]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[16]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[17]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[18]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[19]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[20]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[21]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[22]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[23]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[24]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[25]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[26]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[27]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[28]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[29]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[30]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[31]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[32]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[33]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[34]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[35]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[36]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[37]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[38]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[39]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[40]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[41]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[42]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[43]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[44]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[45]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[46]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[47]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[48]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[49]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[50]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[51]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[52]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[53]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[54]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[55]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[56]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[57]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[58]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[59]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[60]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[61]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[62]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(victimWaymask_lfsr_t[63]); // @[src/main/scala/utils/LFSR64.scala 25:23]
    end
    //
    if (enToggle_past) begin
      cover(io_pf_loadPF_REG_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 284:26]
    end
    //
    if (enToggle_past) begin
      cover(io_pf_storePF_REG_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 285:27]
    end
    //
    if (enToggle_past) begin
      cover(io_pf_laf_REG_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 287:23]
    end
    //
    if (enToggle_past) begin
      cover(io_pf_saf_REG_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 288:23]
    end
    //
    if (enToggle_past) begin
      cover(state_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 298:22]
    end
    //
    if (enToggle_past) begin
      cover(level_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
    end
    //
    if (enToggle_past) begin
      cover(level_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 299:22]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[39]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[40]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[41]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[42]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[43]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[44]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[45]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[46]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[47]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[48]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[49]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[50]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[51]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[52]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[53]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[54]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[55]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[56]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[57]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[58]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[59]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[60]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[61]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[62]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(memRespStore_t[63]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 301:25]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(missMaskStore_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 303:26]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[39]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[40]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[41]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[42]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[43]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[44]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[45]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[46]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[47]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[48]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[49]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[50]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[51]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[52]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[53]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[54]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(raddr_t[55]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 307:18]
    end
    //
    if (enToggle_past) begin
      cover(alreadyOutFire_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 309:33]
    end
    //
    if (enToggle_past) begin
      cover(missPTEAF_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 319:26]
    end
    //
    if (enToggle_past) begin
      cover(REG_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 446:33]
    end
    //
    if (enToggle_past) begin
      cover(REG_1_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:21]
    end
    //
    if (enToggle_past) begin
      cover(REG_1_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:21]
    end
    //
    if (enToggle_past) begin
      cover(REG_1_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:21]
    end
    //
    if (enToggle_past) begin
      cover(REG_1_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:21]
    end
    //
    if (enToggle_past) begin
      cover(REG_2_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:60]
    end
    //
    if (enToggle_past) begin
      cover(REG_2_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:60]
    end
    //
    if (enToggle_past) begin
      cover(REG_2_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:60]
    end
    //
    if (enToggle_past) begin
      cover(REG_2_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:60]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_3_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 447:84]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_4_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_5_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 448:72]
    end
    //
    if (enToggle_past) begin
      cover(REG_6_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_6_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_6_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_6_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_6_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_6_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_6_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_6_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:19]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[39]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[40]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[41]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[42]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_7_t[43]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 449:77]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[39]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[40]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[41]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[42]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[43]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[44]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[45]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[46]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[47]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[48]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[49]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[50]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[51]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[52]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[53]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[54]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(REG_8_t[55]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 450:22]
    end
    //
    if (enToggle_past) begin
      cover(blockRefill_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 453:28]
    end
  end
endmodule
module EmbeddedTLBEmpty_1(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input         io_in_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input  [31:0] io_in_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input  [2:0]  io_in_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input  [3:0]  io_in_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input  [7:0]  io_in_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input  [63:0] io_in_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  input         io_out_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  output        io_out_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  output [2:0]  io_out_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  output [7:0]  io_out_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
  output [63:0] io_out_bits_wdata // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 531:14]
);
  assign io_in_ready = io_out_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
  assign io_out_valid = io_in_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
  assign io_out_bits_addr = io_in_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
  assign io_out_bits_size = io_in_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
  assign io_out_bits_cmd = io_in_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
  assign io_out_bits_wmask = io_in_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
  assign io_out_bits_wdata = io_in_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 536:10]
endmodule
module EmbeddedTLBMD_1(
  input          clock,
  input          reset,
  output [144:0] io_tlbmd_0, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output [144:0] io_tlbmd_1, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output [144:0] io_tlbmd_2, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output [144:0] io_tlbmd_3, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input          io_write_wen, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input  [3:0]   io_write_windex, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input  [3:0]   io_write_waymask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input  [144:0] io_write_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  input  [3:0]   io_rindex, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
  output         io_ready // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 44:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [159:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [144:0] tlbmd_0 [0:15]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_0_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_0_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_0_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_0_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_0_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg [144:0] tlbmd_1 [0:15]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_1_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_1_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_1_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_1_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_1_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg [144:0] tlbmd_2 [0:15]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_2_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_2_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_2_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_2_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_2_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg [144:0] tlbmd_3 [0:15]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_3_MPORT_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_3_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [144:0] tlbmd_3_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire [3:0] tlbmd_3_MPORT_1_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_1_mask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  wire  tlbmd_3_MPORT_1_en; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  reg  resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 56:27]
  reg [3:0] resetSet; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  wrap_wrap = resetSet == 4'hf; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [3:0] _wrap_value_T_1 = resetSet + 4'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  resetFinish = resetState & wrap_wrap; // @[src/main/scala/chisel3/util/Counter.scala 118:{16,23} 117:24]
  wire  _GEN_2 = resetFinish ? 1'h0 : resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 58:22 56:27 58:35]
  wire [3:0] waymask = resetState ? 4'hf : io_write_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 67:20]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  resetState_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 56:27]
  wire  resetState_t = resetState ^ resetState_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 56:27]
  wire  toggle_8065_clock;
  wire  toggle_8065_reset;
  wire  toggle_8065_valid;
  reg  toggle_8065_valid_reg;
  reg [3:0] resetSet_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [3:0] resetSet_t = resetSet ^ resetSet_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  toggle_8066_clock;
  wire  toggle_8066_reset;
  wire [3:0] toggle_8066_valid;
  reg [3:0] toggle_8066_valid_reg;
  GEN_w1_toggle #(.COVER_INDEX(8065)) toggle_8065 (
    .clock(toggle_8065_clock),
    .reset(toggle_8065_reset),
    .valid(toggle_8065_valid)
  );
  GEN_w4_toggle #(.COVER_INDEX(8066)) toggle_8066 (
    .clock(toggle_8066_clock),
    .reset(toggle_8066_reset),
    .valid(toggle_8066_valid)
  );
  assign tlbmd_0_MPORT_en = 1'h1;
  assign tlbmd_0_MPORT_addr = io_rindex;
  assign tlbmd_0_MPORT_data = tlbmd_0[tlbmd_0_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_0_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_0_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_0_MPORT_1_mask = waymask[0];
  assign tlbmd_0_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_1_MPORT_en = 1'h1;
  assign tlbmd_1_MPORT_addr = io_rindex;
  assign tlbmd_1_MPORT_data = tlbmd_1[tlbmd_1_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_1_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_1_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_1_MPORT_1_mask = waymask[1];
  assign tlbmd_1_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_2_MPORT_en = 1'h1;
  assign tlbmd_2_MPORT_addr = io_rindex;
  assign tlbmd_2_MPORT_data = tlbmd_2[tlbmd_2_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_2_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_2_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_2_MPORT_1_mask = waymask[2];
  assign tlbmd_2_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_3_MPORT_en = 1'h1;
  assign tlbmd_3_MPORT_addr = io_rindex;
  assign tlbmd_3_MPORT_data = tlbmd_3[tlbmd_3_MPORT_addr]; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
  assign tlbmd_3_MPORT_1_data = resetState ? 145'h0 : io_write_wdata;
  assign tlbmd_3_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_3_MPORT_1_mask = waymask[3];
  assign tlbmd_3_MPORT_1_en = resetState | io_write_wen;
  assign io_tlbmd_0 = tlbmd_0_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_tlbmd_1 = tlbmd_1_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_tlbmd_2 = tlbmd_2_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_tlbmd_3 = tlbmd_3_MPORT_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 53:12]
  assign io_ready = ~resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 73:15]
  assign toggle_8065_clock = clock;
  assign toggle_8065_reset = reset;
  assign toggle_8065_valid = resetState ^ toggle_8065_valid_reg;
  assign toggle_8066_clock = clock;
  assign toggle_8066_reset = reset;
  assign toggle_8066_valid = resetSet ^ toggle_8066_valid_reg;
  always @(posedge clock) begin
    if (tlbmd_0_MPORT_1_en & tlbmd_0_MPORT_1_mask) begin
      tlbmd_0[tlbmd_0_MPORT_1_addr] <= tlbmd_0_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    if (tlbmd_1_MPORT_1_en & tlbmd_1_MPORT_1_mask) begin
      tlbmd_1[tlbmd_1_MPORT_1_addr] <= tlbmd_1_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    if (tlbmd_2_MPORT_1_en & tlbmd_2_MPORT_1_mask) begin
      tlbmd_2[tlbmd_2_MPORT_1_addr] <= tlbmd_2_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    if (tlbmd_3_MPORT_1_en & tlbmd_3_MPORT_1_mask) begin
      tlbmd_3[tlbmd_3_MPORT_1_addr] <= tlbmd_3_MPORT_1_data; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 52:18]
    end
    resetState <= reset | _GEN_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 56:{27,27}]
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      resetSet <= 4'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (resetState) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      resetSet <= _wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    resetState_p <= resetState; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 56:27]
    toggle_8065_valid_reg <= resetState;
    resetSet_p <= resetSet; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    toggle_8066_valid_reg <= resetSet;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {5{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_0[initvar] = _RAND_0[144:0];
  _RAND_1 = {5{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_1[initvar] = _RAND_1[144:0];
  _RAND_2 = {5{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_2[initvar] = _RAND_2[144:0];
  _RAND_3 = {5{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_3[initvar] = _RAND_3[144:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  resetState = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  resetSet = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  resetState_p = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  toggle_8065_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  resetSet_p = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  toggle_8066_valid_reg = _RAND_9[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(resetState_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 56:27]
    end
    //
    if (enToggle_past) begin
      cover(resetSet_t[0]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(resetSet_t[1]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(resetSet_t[2]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(resetSet_t[3]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
  end
endmodule
module EmbeddedTLB_1(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [38:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [2:0]  io_in_req_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_out_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_out_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [2:0]  io_out_req_bits_size, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_out_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [63:0] io_out_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_mem_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_mem_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [31:0] io_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [3:0]  io_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output [63:0] io_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_mem_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [63:0] io_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input  [1:0]  io_csrMMU_priviledgeMode, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_csrMMU_status_sum, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         io_csrMMU_status_mxr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_csrMMU_loadPF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_csrMMU_storePF, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_csrMMU_laf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  output        io_csrMMU_saf, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 40:14]
  input         lr,
  input         scInflight,
  input         amoReq,
  input  [63:0] lrAddr,
  output [55:0] paddr,
  input  [63:0] CSRSATP,
  output        _T_12_0,
  output        scIsSuccess_0,
  output        vmEnable_0,
  input         MOUFlushTLB,
  output        tlbFinish_0,
  output        _T_13_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [159:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [159:0] _RAND_17;
  reg [159:0] _RAND_18;
  reg [159:0] _RAND_19;
  reg [159:0] _RAND_20;
  reg [159:0] _RAND_21;
  reg [159:0] _RAND_22;
  reg [159:0] _RAND_23;
  reg [159:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
`endif // RANDOMIZE_REG_INIT
  wire  tlbExec_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_in_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [38:0] tlbExec_io_in_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [2:0] tlbExec_io_in_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_in_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [7:0] tlbExec_io_in_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_in_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_out_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_out_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [31:0] tlbExec_io_out_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [2:0] tlbExec_io_out_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [7:0] tlbExec_io_out_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_out_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_md_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mdWrite_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_mdWrite_windex; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_mdWrite_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [144:0] tlbExec_io_mdWrite_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mdReady; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [31:0] tlbExec_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [3:0] tlbExec_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_io_satp; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [1:0] tlbExec_io_pf_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_status_sum; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_status_mxr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_laf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_pf_saf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_io_isFinish; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_lr_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_scInflight_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_ISAMO; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [63:0] tlbExec_lr_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire [55:0] tlbExec_paddr_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbExec_scIsSuccess_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
  wire  tlbEmpty_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire  tlbEmpty_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire  tlbEmpty_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire  tlbEmpty_io_in_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [31:0] tlbEmpty_io_in_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [2:0] tlbEmpty_io_in_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [3:0] tlbEmpty_io_in_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [7:0] tlbEmpty_io_in_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [63:0] tlbEmpty_io_in_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire  tlbEmpty_io_out_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire  tlbEmpty_io_out_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [31:0] tlbEmpty_io_out_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [2:0] tlbEmpty_io_out_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [3:0] tlbEmpty_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [7:0] tlbEmpty_io_out_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire [63:0] tlbEmpty_io_out_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
  wire  mdTLB_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  mdTLB_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_tlbmd_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  mdTLB_io_write_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [3:0] mdTLB_io_write_windex; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [3:0] mdTLB_io_write_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [144:0] mdTLB_io_write_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire [3:0] mdTLB_io_rindex; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  mdTLB_io_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
  wire  vmEnable = CSRSATP[63:60] == 4'h8 & io_csrMMU_priviledgeMode < 2'h3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 90:57]
  reg [144:0] r_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  reg [144:0] r_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  reg [144:0] r_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  reg [144:0] r_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire  mdUpdate = io_in_req_valid & tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 116:26]
  reg  valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
  wire  _GEN_7 = tlbExec_io_isFinish ? 1'h0 : valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24 108:{25,33}]
  wire  _GEN_8 = mdUpdate & vmEnable | _GEN_7; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 109:{50,58}]
  reg [38:0] tlbExec_io_in_bits_r_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  reg [2:0] tlbExec_io_in_bits_r_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  reg [3:0] tlbExec_io_in_bits_r_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  reg [7:0] tlbExec_io_in_bits_r_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  reg [63:0] tlbExec_io_in_bits_r_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  wire  _T_7 = tlbEmpty_io_out_ready & tlbEmpty_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  _GEN_15 = _T_7 ? 1'h0 : valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24 25:{25,33}]
  wire  _T_8 = tlbExec_io_out_valid & tlbEmpty_io_in_ready; // @[src/main/scala/utils/Pipeline.scala 26:22]
  wire  _GEN_16 = tlbExec_io_out_valid & tlbEmpty_io_in_ready | _GEN_15; // @[src/main/scala/utils/Pipeline.scala 26:{38,46}]
  reg [31:0] tlbEmpty_io_in_bits_r_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [2:0] tlbEmpty_io_in_bits_r_size; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [3:0] tlbEmpty_io_in_bits_r_cmd; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [7:0] tlbEmpty_io_in_bits_r_wmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg [63:0] tlbEmpty_io_in_bits_r_wdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
  reg  alreadyOutFinish; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 176:37]
  wire  _GEN_36 = tlbExec_io_out_valid & ~tlbExec_io_out_ready | alreadyOutFinish; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 176:{37,37,37}]
  wire  _T_10 = tlbExec_io_out_ready & tlbExec_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _tlbFinish_T_2 = tlbExec_io_pf_loadPF | tlbExec_io_pf_storePF; // @[src/main/scala/nutcore/Bundle.scala 134:23]
  wire  _tlbFinish_T_3 = tlbExec_io_pf_laf | tlbExec_io_pf_saf; // @[src/main/scala/nutcore/Bundle.scala 135:24]
  wire  _tlbFinish_T_4 = _tlbFinish_T_2 | _tlbFinish_T_3; // @[src/main/scala/nutcore/Bundle.scala 136:35]
  wire  tlbFinish = tlbExec_io_out_valid & ~alreadyOutFinish | _tlbFinish_T_4 | ~scIsSuccess_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 180:95]
  wire  _T_12 = io_csrMMU_loadPF | io_csrMMU_storePF; // @[src/main/scala/nutcore/Bundle.scala 134:23]
  wire  _T_13 = io_csrMMU_laf | io_csrMMU_saf; // @[src/main/scala/nutcore/Bundle.scala 135:24]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [144:0] r_0_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire [144:0] r_0_t = r_0 ^ r_0_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire  toggle_8070_clock;
  wire  toggle_8070_reset;
  wire [144:0] toggle_8070_valid;
  reg [144:0] toggle_8070_valid_reg;
  reg [144:0] r_1_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire [144:0] r_1_t = r_1 ^ r_1_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire  toggle_8215_clock;
  wire  toggle_8215_reset;
  wire [144:0] toggle_8215_valid;
  reg [144:0] toggle_8215_valid_reg;
  reg [144:0] r_2_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire [144:0] r_2_t = r_2 ^ r_2_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire  toggle_8360_clock;
  wire  toggle_8360_reset;
  wire [144:0] toggle_8360_valid;
  reg [144:0] toggle_8360_valid_reg;
  reg [144:0] r_3_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire [144:0] r_3_t = r_3 ^ r_3_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
  wire  toggle_8505_clock;
  wire  toggle_8505_reset;
  wire [144:0] toggle_8505_valid;
  reg [144:0] toggle_8505_valid_reg;
  reg  valid_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
  wire  valid_t = valid ^ valid_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
  wire  toggle_8650_clock;
  wire  toggle_8650_reset;
  wire  toggle_8650_valid;
  reg  toggle_8650_valid_reg;
  reg [38:0] tlbExec_io_in_bits_r_addr_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  wire [38:0] tlbExec_io_in_bits_r_addr_t = tlbExec_io_in_bits_r_addr ^ tlbExec_io_in_bits_r_addr_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  wire  toggle_8651_clock;
  wire  toggle_8651_reset;
  wire [38:0] toggle_8651_valid;
  reg [38:0] toggle_8651_valid_reg;
  reg [2:0] tlbExec_io_in_bits_r_size_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  wire [2:0] tlbExec_io_in_bits_r_size_t = tlbExec_io_in_bits_r_size ^ tlbExec_io_in_bits_r_size_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  wire  toggle_8690_clock;
  wire  toggle_8690_reset;
  wire [2:0] toggle_8690_valid;
  reg [2:0] toggle_8690_valid_reg;
  reg [3:0] tlbExec_io_in_bits_r_cmd_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  wire [3:0] tlbExec_io_in_bits_r_cmd_t = tlbExec_io_in_bits_r_cmd ^ tlbExec_io_in_bits_r_cmd_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  wire  toggle_8693_clock;
  wire  toggle_8693_reset;
  wire [3:0] toggle_8693_valid;
  reg [3:0] toggle_8693_valid_reg;
  reg [7:0] tlbExec_io_in_bits_r_wmask_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  wire [7:0] tlbExec_io_in_bits_r_wmask_t = tlbExec_io_in_bits_r_wmask ^ tlbExec_io_in_bits_r_wmask_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  wire  toggle_8697_clock;
  wire  toggle_8697_reset;
  wire [7:0] toggle_8697_valid;
  reg [7:0] toggle_8697_valid_reg;
  reg [63:0] tlbExec_io_in_bits_r_wdata_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  wire [63:0] tlbExec_io_in_bits_r_wdata_t = tlbExec_io_in_bits_r_wdata ^ tlbExec_io_in_bits_r_wdata_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
  wire  toggle_8705_clock;
  wire  toggle_8705_reset;
  wire [63:0] toggle_8705_valid;
  reg [63:0] toggle_8705_valid_reg;
  reg  valid_1_p; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  valid_1_t = valid_1 ^ valid_1_p; // @[src/main/scala/utils/Pipeline.scala 24:24]
  wire  toggle_8769_clock;
  wire  toggle_8769_reset;
  wire  toggle_8769_valid;
  reg  toggle_8769_valid_reg;
  reg [31:0] tlbEmpty_io_in_bits_r_addr_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [31:0] tlbEmpty_io_in_bits_r_addr_t = tlbEmpty_io_in_bits_r_addr ^ tlbEmpty_io_in_bits_r_addr_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_8770_clock;
  wire  toggle_8770_reset;
  wire [31:0] toggle_8770_valid;
  reg [31:0] toggle_8770_valid_reg;
  reg [2:0] tlbEmpty_io_in_bits_r_size_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [2:0] tlbEmpty_io_in_bits_r_size_t = tlbEmpty_io_in_bits_r_size ^ tlbEmpty_io_in_bits_r_size_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_8802_clock;
  wire  toggle_8802_reset;
  wire [2:0] toggle_8802_valid;
  reg [2:0] toggle_8802_valid_reg;
  reg [3:0] tlbEmpty_io_in_bits_r_cmd_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [3:0] tlbEmpty_io_in_bits_r_cmd_t = tlbEmpty_io_in_bits_r_cmd ^ tlbEmpty_io_in_bits_r_cmd_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_8805_clock;
  wire  toggle_8805_reset;
  wire [3:0] toggle_8805_valid;
  reg [3:0] toggle_8805_valid_reg;
  reg [7:0] tlbEmpty_io_in_bits_r_wmask_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [7:0] tlbEmpty_io_in_bits_r_wmask_t = tlbEmpty_io_in_bits_r_wmask ^ tlbEmpty_io_in_bits_r_wmask_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_8809_clock;
  wire  toggle_8809_reset;
  wire [7:0] toggle_8809_valid;
  reg [7:0] toggle_8809_valid_reg;
  reg [63:0] tlbEmpty_io_in_bits_r_wdata_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire [63:0] tlbEmpty_io_in_bits_r_wdata_t = tlbEmpty_io_in_bits_r_wdata ^ tlbEmpty_io_in_bits_r_wdata_p; // @[src/main/scala/utils/Pipeline.scala 30:28]
  wire  toggle_8817_clock;
  wire  toggle_8817_reset;
  wire [63:0] toggle_8817_valid;
  reg [63:0] toggle_8817_valid_reg;
  reg  alreadyOutFinish_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 176:37]
  wire  alreadyOutFinish_t = alreadyOutFinish ^ alreadyOutFinish_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 176:37]
  wire  toggle_8881_clock;
  wire  toggle_8881_reset;
  wire  toggle_8881_valid;
  reg  toggle_8881_valid_reg;
  EmbeddedTLBExec_1 tlbExec ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 84:23]
    .clock(tlbExec_clock),
    .reset(tlbExec_reset),
    .io_in_ready(tlbExec_io_in_ready),
    .io_in_valid(tlbExec_io_in_valid),
    .io_in_bits_addr(tlbExec_io_in_bits_addr),
    .io_in_bits_size(tlbExec_io_in_bits_size),
    .io_in_bits_cmd(tlbExec_io_in_bits_cmd),
    .io_in_bits_wmask(tlbExec_io_in_bits_wmask),
    .io_in_bits_wdata(tlbExec_io_in_bits_wdata),
    .io_out_ready(tlbExec_io_out_ready),
    .io_out_valid(tlbExec_io_out_valid),
    .io_out_bits_addr(tlbExec_io_out_bits_addr),
    .io_out_bits_size(tlbExec_io_out_bits_size),
    .io_out_bits_cmd(tlbExec_io_out_bits_cmd),
    .io_out_bits_wmask(tlbExec_io_out_bits_wmask),
    .io_out_bits_wdata(tlbExec_io_out_bits_wdata),
    .io_md_0(tlbExec_io_md_0),
    .io_md_1(tlbExec_io_md_1),
    .io_md_2(tlbExec_io_md_2),
    .io_md_3(tlbExec_io_md_3),
    .io_mdWrite_wen(tlbExec_io_mdWrite_wen),
    .io_mdWrite_windex(tlbExec_io_mdWrite_windex),
    .io_mdWrite_waymask(tlbExec_io_mdWrite_waymask),
    .io_mdWrite_wdata(tlbExec_io_mdWrite_wdata),
    .io_mdReady(tlbExec_io_mdReady),
    .io_mem_req_ready(tlbExec_io_mem_req_ready),
    .io_mem_req_valid(tlbExec_io_mem_req_valid),
    .io_mem_req_bits_addr(tlbExec_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(tlbExec_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(tlbExec_io_mem_req_bits_wdata),
    .io_mem_resp_ready(tlbExec_io_mem_resp_ready),
    .io_mem_resp_valid(tlbExec_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(tlbExec_io_mem_resp_bits_rdata),
    .io_satp(tlbExec_io_satp),
    .io_pf_priviledgeMode(tlbExec_io_pf_priviledgeMode),
    .io_pf_status_sum(tlbExec_io_pf_status_sum),
    .io_pf_status_mxr(tlbExec_io_pf_status_mxr),
    .io_pf_loadPF(tlbExec_io_pf_loadPF),
    .io_pf_storePF(tlbExec_io_pf_storePF),
    .io_pf_laf(tlbExec_io_pf_laf),
    .io_pf_saf(tlbExec_io_pf_saf),
    .io_isFinish(tlbExec_io_isFinish),
    .lr_0(tlbExec_lr_0),
    .scInflight_0(tlbExec_scInflight_0),
    .ISAMO(tlbExec_ISAMO),
    .lr_addr(tlbExec_lr_addr),
    .paddr_0(tlbExec_paddr_0),
    .scIsSuccess_0(tlbExec_scIsSuccess_0)
  );
  EmbeddedTLBEmpty_1 tlbEmpty ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 85:24]
    .clock(tlbEmpty_clock),
    .reset(tlbEmpty_reset),
    .io_in_ready(tlbEmpty_io_in_ready),
    .io_in_valid(tlbEmpty_io_in_valid),
    .io_in_bits_addr(tlbEmpty_io_in_bits_addr),
    .io_in_bits_size(tlbEmpty_io_in_bits_size),
    .io_in_bits_cmd(tlbEmpty_io_in_bits_cmd),
    .io_in_bits_wmask(tlbEmpty_io_in_bits_wmask),
    .io_in_bits_wdata(tlbEmpty_io_in_bits_wdata),
    .io_out_ready(tlbEmpty_io_out_ready),
    .io_out_valid(tlbEmpty_io_out_valid),
    .io_out_bits_addr(tlbEmpty_io_out_bits_addr),
    .io_out_bits_size(tlbEmpty_io_out_bits_size),
    .io_out_bits_cmd(tlbEmpty_io_out_bits_cmd),
    .io_out_bits_wmask(tlbEmpty_io_out_bits_wmask),
    .io_out_bits_wdata(tlbEmpty_io_out_bits_wdata)
  );
  EmbeddedTLBMD_1 mdTLB ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 86:21]
    .clock(mdTLB_clock),
    .reset(mdTLB_reset),
    .io_tlbmd_0(mdTLB_io_tlbmd_0),
    .io_tlbmd_1(mdTLB_io_tlbmd_1),
    .io_tlbmd_2(mdTLB_io_tlbmd_2),
    .io_tlbmd_3(mdTLB_io_tlbmd_3),
    .io_write_wen(mdTLB_io_write_wen),
    .io_write_windex(mdTLB_io_write_windex),
    .io_write_waymask(mdTLB_io_write_waymask),
    .io_write_wdata(mdTLB_io_write_wdata),
    .io_rindex(mdTLB_io_rindex),
    .io_ready(mdTLB_io_ready)
  );
  GEN_w145_toggle #(.COVER_INDEX(8070)) toggle_8070 (
    .clock(toggle_8070_clock),
    .reset(toggle_8070_reset),
    .valid(toggle_8070_valid)
  );
  GEN_w145_toggle #(.COVER_INDEX(8215)) toggle_8215 (
    .clock(toggle_8215_clock),
    .reset(toggle_8215_reset),
    .valid(toggle_8215_valid)
  );
  GEN_w145_toggle #(.COVER_INDEX(8360)) toggle_8360 (
    .clock(toggle_8360_clock),
    .reset(toggle_8360_reset),
    .valid(toggle_8360_valid)
  );
  GEN_w145_toggle #(.COVER_INDEX(8505)) toggle_8505 (
    .clock(toggle_8505_clock),
    .reset(toggle_8505_reset),
    .valid(toggle_8505_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(8650)) toggle_8650 (
    .clock(toggle_8650_clock),
    .reset(toggle_8650_reset),
    .valid(toggle_8650_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(8651)) toggle_8651 (
    .clock(toggle_8651_clock),
    .reset(toggle_8651_reset),
    .valid(toggle_8651_valid)
  );
  GEN_w3_toggle #(.COVER_INDEX(8690)) toggle_8690 (
    .clock(toggle_8690_clock),
    .reset(toggle_8690_reset),
    .valid(toggle_8690_valid)
  );
  GEN_w4_toggle #(.COVER_INDEX(8693)) toggle_8693 (
    .clock(toggle_8693_clock),
    .reset(toggle_8693_reset),
    .valid(toggle_8693_valid)
  );
  GEN_w8_toggle #(.COVER_INDEX(8697)) toggle_8697 (
    .clock(toggle_8697_clock),
    .reset(toggle_8697_reset),
    .valid(toggle_8697_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(8705)) toggle_8705 (
    .clock(toggle_8705_clock),
    .reset(toggle_8705_reset),
    .valid(toggle_8705_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(8769)) toggle_8769 (
    .clock(toggle_8769_clock),
    .reset(toggle_8769_reset),
    .valid(toggle_8769_valid)
  );
  GEN_w32_toggle #(.COVER_INDEX(8770)) toggle_8770 (
    .clock(toggle_8770_clock),
    .reset(toggle_8770_reset),
    .valid(toggle_8770_valid)
  );
  GEN_w3_toggle #(.COVER_INDEX(8802)) toggle_8802 (
    .clock(toggle_8802_clock),
    .reset(toggle_8802_reset),
    .valid(toggle_8802_valid)
  );
  GEN_w4_toggle #(.COVER_INDEX(8805)) toggle_8805 (
    .clock(toggle_8805_clock),
    .reset(toggle_8805_reset),
    .valid(toggle_8805_valid)
  );
  GEN_w8_toggle #(.COVER_INDEX(8809)) toggle_8809 (
    .clock(toggle_8809_clock),
    .reset(toggle_8809_reset),
    .valid(toggle_8809_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(8817)) toggle_8817 (
    .clock(toggle_8817_clock),
    .reset(toggle_8817_reset),
    .valid(toggle_8817_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(8881)) toggle_8881 (
    .clock(toggle_8881_clock),
    .reset(toggle_8881_reset),
    .valid(toggle_8881_valid)
  );
  assign io_in_req_ready = ~vmEnable ? io_out_req_ready : tlbExec_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 112:16 144:19 149:23]
  assign io_in_resp_valid = io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 172:15]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 172:15]
  assign io_out_req_valid = ~vmEnable ? io_in_req_valid : tlbEmpty_io_out_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 148:24 169:41]
  assign io_out_req_bits_addr = ~vmEnable ? io_in_req_bits_addr[31:0] : tlbEmpty_io_out_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 162:26 169:41]
  assign io_out_req_bits_size = ~vmEnable ? io_in_req_bits_size : tlbEmpty_io_out_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 163:26 169:41]
  assign io_out_req_bits_cmd = ~vmEnable ? io_in_req_bits_cmd : tlbEmpty_io_out_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 164:25 169:41]
  assign io_out_req_bits_wmask = ~vmEnable ? io_in_req_bits_wmask : tlbEmpty_io_out_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 165:27 169:41]
  assign io_out_req_bits_wdata = ~vmEnable ? io_in_req_bits_wdata : tlbEmpty_io_out_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 166:27 169:41]
  assign io_mem_req_valid = tlbExec_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_mem_req_bits_addr = tlbExec_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_mem_req_bits_cmd = tlbExec_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_mem_req_bits_wdata = tlbExec_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign io_csrMMU_loadPF = ~vmEnable ? 1'h0 : tlbExec_io_pf_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 150:24 95:17]
  assign io_csrMMU_storePF = ~vmEnable ? 1'h0 : tlbExec_io_pf_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 151:25 95:17]
  assign io_csrMMU_laf = ~vmEnable ? 1'h0 : tlbExec_io_pf_laf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 152:21 95:17]
  assign io_csrMMU_saf = ~vmEnable ? 1'h0 : tlbExec_io_pf_saf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 153:21 95:17]
  assign paddr = tlbExec_paddr_0;
  assign _T_12_0 = _T_12;
  assign scIsSuccess_0 = tlbExec_scIsSuccess_0;
  assign vmEnable_0 = vmEnable;
  assign tlbFinish_0 = tlbFinish;
  assign _T_13_1 = _T_13;
  assign tlbExec_clock = clock;
  assign tlbExec_reset = reset;
  assign tlbExec_io_in_valid = valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 114:17]
  assign tlbExec_io_in_bits_addr = tlbExec_io_in_bits_r_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_in_bits_size = tlbExec_io_in_bits_r_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_in_bits_cmd = tlbExec_io_in_bits_r_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_in_bits_wmask = tlbExec_io_in_bits_r_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_in_bits_wdata = tlbExec_io_in_bits_r_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:16]
  assign tlbExec_io_out_ready = ~vmEnable | tlbEmpty_io_in_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 145:26 src/main/scala/utils/Pipeline.scala 29:16]
  assign tlbExec_io_md_0 = r_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_md_1 = r_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_md_2 = r_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_md_3 = r_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:17]
  assign tlbExec_io_mdReady = mdTLB_io_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 97:22]
  assign tlbExec_io_mem_req_ready = io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign tlbExec_io_mem_resp_valid = io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign tlbExec_io_mem_resp_bits_rdata = io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 94:18]
  assign tlbExec_io_satp = CSRSATP; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 80:22]
  assign tlbExec_io_pf_priviledgeMode = io_csrMMU_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 95:17]
  assign tlbExec_io_pf_status_sum = io_csrMMU_status_sum; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 95:17]
  assign tlbExec_io_pf_status_mxr = io_csrMMU_status_mxr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 95:17]
  assign tlbExec_lr_0 = lr;
  assign tlbExec_scInflight_0 = scInflight;
  assign tlbExec_ISAMO = amoReq;
  assign tlbExec_lr_addr = lrAddr;
  assign tlbEmpty_clock = clock;
  assign tlbEmpty_reset = reset;
  assign tlbEmpty_io_in_valid = valid_1; // @[src/main/scala/utils/Pipeline.scala 31:17]
  assign tlbEmpty_io_in_bits_addr = tlbEmpty_io_in_bits_r_addr; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_size = tlbEmpty_io_in_bits_r_size; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_cmd = tlbEmpty_io_in_bits_r_cmd; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_wmask = tlbEmpty_io_in_bits_r_wmask; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_wdata = tlbEmpty_io_in_bits_r_wdata; // @[src/main/scala/utils/Pipeline.scala 30:16]
  assign tlbEmpty_io_out_ready = ~vmEnable | io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 144:19 147:29 169:41]
  assign mdTLB_clock = clock;
  assign mdTLB_reset = reset | MOUFlushTLB; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 104:31]
  assign mdTLB_io_write_wen = tlbExec_io_mdWrite_wen; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  assign mdTLB_io_write_windex = tlbExec_io_mdWrite_windex; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  assign mdTLB_io_write_waymask = tlbExec_io_mdWrite_waymask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  assign mdTLB_io_write_wdata = tlbExec_io_mdWrite_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 99:18]
  assign mdTLB_io_rindex = io_in_req_bits_addr[15:12]; // @[src/main/scala/nutcore/mem/TLB.scala 203:19]
  assign toggle_8070_clock = clock;
  assign toggle_8070_reset = reset;
  assign toggle_8070_valid = r_0 ^ toggle_8070_valid_reg;
  assign toggle_8215_clock = clock;
  assign toggle_8215_reset = reset;
  assign toggle_8215_valid = r_1 ^ toggle_8215_valid_reg;
  assign toggle_8360_clock = clock;
  assign toggle_8360_reset = reset;
  assign toggle_8360_valid = r_2 ^ toggle_8360_valid_reg;
  assign toggle_8505_clock = clock;
  assign toggle_8505_reset = reset;
  assign toggle_8505_valid = r_3 ^ toggle_8505_valid_reg;
  assign toggle_8650_clock = clock;
  assign toggle_8650_reset = reset;
  assign toggle_8650_valid = valid ^ toggle_8650_valid_reg;
  assign toggle_8651_clock = clock;
  assign toggle_8651_reset = reset;
  assign toggle_8651_valid = tlbExec_io_in_bits_r_addr ^ toggle_8651_valid_reg;
  assign toggle_8690_clock = clock;
  assign toggle_8690_reset = reset;
  assign toggle_8690_valid = tlbExec_io_in_bits_r_size ^ toggle_8690_valid_reg;
  assign toggle_8693_clock = clock;
  assign toggle_8693_reset = reset;
  assign toggle_8693_valid = tlbExec_io_in_bits_r_cmd ^ toggle_8693_valid_reg;
  assign toggle_8697_clock = clock;
  assign toggle_8697_reset = reset;
  assign toggle_8697_valid = tlbExec_io_in_bits_r_wmask ^ toggle_8697_valid_reg;
  assign toggle_8705_clock = clock;
  assign toggle_8705_reset = reset;
  assign toggle_8705_valid = tlbExec_io_in_bits_r_wdata ^ toggle_8705_valid_reg;
  assign toggle_8769_clock = clock;
  assign toggle_8769_reset = reset;
  assign toggle_8769_valid = valid_1 ^ toggle_8769_valid_reg;
  assign toggle_8770_clock = clock;
  assign toggle_8770_reset = reset;
  assign toggle_8770_valid = tlbEmpty_io_in_bits_r_addr ^ toggle_8770_valid_reg;
  assign toggle_8802_clock = clock;
  assign toggle_8802_reset = reset;
  assign toggle_8802_valid = tlbEmpty_io_in_bits_r_size ^ toggle_8802_valid_reg;
  assign toggle_8805_clock = clock;
  assign toggle_8805_reset = reset;
  assign toggle_8805_valid = tlbEmpty_io_in_bits_r_cmd ^ toggle_8805_valid_reg;
  assign toggle_8809_clock = clock;
  assign toggle_8809_reset = reset;
  assign toggle_8809_valid = tlbEmpty_io_in_bits_r_wmask ^ toggle_8809_valid_reg;
  assign toggle_8817_clock = clock;
  assign toggle_8817_reset = reset;
  assign toggle_8817_valid = tlbEmpty_io_in_bits_r_wdata ^ toggle_8817_valid_reg;
  assign toggle_8881_clock = clock;
  assign toggle_8881_reset = reset;
  assign toggle_8881_valid = alreadyOutFinish ^ toggle_8881_valid_reg;
  always @(posedge clock) begin
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_0 <= mdTLB_io_tlbmd_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_1 <= mdTLB_io_tlbmd_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_2 <= mdTLB_io_tlbmd_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
      r_3 <= mdTLB_io_tlbmd_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
      valid <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
    end else begin
      valid <= _GEN_8;
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_addr <= io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_size <= io_in_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_cmd <= io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_wmask <= io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    if (mdUpdate) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
      tlbExec_io_in_bits_r_wdata <= io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    if (reset) begin // @[src/main/scala/utils/Pipeline.scala 24:24]
      valid_1 <= 1'h0; // @[src/main/scala/utils/Pipeline.scala 24:24]
    end else begin
      valid_1 <= _GEN_16;
    end
    if (_T_8) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      tlbEmpty_io_in_bits_r_addr <= tlbExec_io_out_bits_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_8) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      tlbEmpty_io_in_bits_r_size <= tlbExec_io_out_bits_size; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_8) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      tlbEmpty_io_in_bits_r_cmd <= tlbExec_io_out_bits_cmd; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_8) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      tlbEmpty_io_in_bits_r_wmask <= tlbExec_io_out_bits_wmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (_T_8) begin // @[src/main/scala/utils/Pipeline.scala 30:28]
      tlbEmpty_io_in_bits_r_wdata <= tlbExec_io_out_bits_wdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 176:37]
      alreadyOutFinish <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 176:37]
    end else if (alreadyOutFinish & _T_10) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 177:53]
      alreadyOutFinish <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 177:72]
    end else begin
      alreadyOutFinish <= _GEN_36;
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    r_0_p <= r_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    toggle_8070_valid_reg <= r_0;
    r_1_p <= r_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    toggle_8215_valid_reg <= r_1;
    r_2_p <= r_2; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    toggle_8360_valid_reg <= r_2;
    r_3_p <= r_3; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    toggle_8505_valid_reg <= r_3;
    valid_p <= valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
    toggle_8650_valid_reg <= valid;
    tlbExec_io_in_bits_r_addr_p <= tlbExec_io_in_bits_r_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    toggle_8651_valid_reg <= tlbExec_io_in_bits_r_addr;
    tlbExec_io_in_bits_r_size_p <= tlbExec_io_in_bits_r_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    toggle_8690_valid_reg <= tlbExec_io_in_bits_r_size;
    tlbExec_io_in_bits_r_cmd_p <= tlbExec_io_in_bits_r_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    toggle_8693_valid_reg <= tlbExec_io_in_bits_r_cmd;
    tlbExec_io_in_bits_r_wmask_p <= tlbExec_io_in_bits_r_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    toggle_8697_valid_reg <= tlbExec_io_in_bits_r_wmask;
    tlbExec_io_in_bits_r_wdata_p <= tlbExec_io_in_bits_r_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    toggle_8705_valid_reg <= tlbExec_io_in_bits_r_wdata;
    valid_1_p <= valid_1; // @[src/main/scala/utils/Pipeline.scala 24:24]
    toggle_8769_valid_reg <= valid_1;
    tlbEmpty_io_in_bits_r_addr_p <= tlbEmpty_io_in_bits_r_addr; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_8770_valid_reg <= tlbEmpty_io_in_bits_r_addr;
    tlbEmpty_io_in_bits_r_size_p <= tlbEmpty_io_in_bits_r_size; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_8802_valid_reg <= tlbEmpty_io_in_bits_r_size;
    tlbEmpty_io_in_bits_r_cmd_p <= tlbEmpty_io_in_bits_r_cmd; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_8805_valid_reg <= tlbEmpty_io_in_bits_r_cmd;
    tlbEmpty_io_in_bits_r_wmask_p <= tlbEmpty_io_in_bits_r_wmask; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_8809_valid_reg <= tlbEmpty_io_in_bits_r_wmask;
    tlbEmpty_io_in_bits_r_wdata_p <= tlbEmpty_io_in_bits_r_wdata; // @[src/main/scala/utils/Pipeline.scala 30:28]
    toggle_8817_valid_reg <= tlbEmpty_io_in_bits_r_wdata;
    alreadyOutFinish_p <= alreadyOutFinish; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 176:37]
    toggle_8881_valid_reg <= alreadyOutFinish;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {5{`RANDOM}};
  r_0 = _RAND_0[144:0];
  _RAND_1 = {5{`RANDOM}};
  r_1 = _RAND_1[144:0];
  _RAND_2 = {5{`RANDOM}};
  r_2 = _RAND_2[144:0];
  _RAND_3 = {5{`RANDOM}};
  r_3 = _RAND_3[144:0];
  _RAND_4 = {1{`RANDOM}};
  valid = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  tlbExec_io_in_bits_r_addr = _RAND_5[38:0];
  _RAND_6 = {1{`RANDOM}};
  tlbExec_io_in_bits_r_size = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  tlbExec_io_in_bits_r_cmd = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  tlbExec_io_in_bits_r_wmask = _RAND_8[7:0];
  _RAND_9 = {2{`RANDOM}};
  tlbExec_io_in_bits_r_wdata = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  valid_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  tlbEmpty_io_in_bits_r_addr = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  tlbEmpty_io_in_bits_r_size = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  tlbEmpty_io_in_bits_r_cmd = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  tlbEmpty_io_in_bits_r_wmask = _RAND_14[7:0];
  _RAND_15 = {2{`RANDOM}};
  tlbEmpty_io_in_bits_r_wdata = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  alreadyOutFinish = _RAND_16[0:0];
  _RAND_17 = {5{`RANDOM}};
  r_0_p = _RAND_17[144:0];
  _RAND_18 = {5{`RANDOM}};
  toggle_8070_valid_reg = _RAND_18[144:0];
  _RAND_19 = {5{`RANDOM}};
  r_1_p = _RAND_19[144:0];
  _RAND_20 = {5{`RANDOM}};
  toggle_8215_valid_reg = _RAND_20[144:0];
  _RAND_21 = {5{`RANDOM}};
  r_2_p = _RAND_21[144:0];
  _RAND_22 = {5{`RANDOM}};
  toggle_8360_valid_reg = _RAND_22[144:0];
  _RAND_23 = {5{`RANDOM}};
  r_3_p = _RAND_23[144:0];
  _RAND_24 = {5{`RANDOM}};
  toggle_8505_valid_reg = _RAND_24[144:0];
  _RAND_25 = {1{`RANDOM}};
  valid_p = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  toggle_8650_valid_reg = _RAND_26[0:0];
  _RAND_27 = {2{`RANDOM}};
  tlbExec_io_in_bits_r_addr_p = _RAND_27[38:0];
  _RAND_28 = {2{`RANDOM}};
  toggle_8651_valid_reg = _RAND_28[38:0];
  _RAND_29 = {1{`RANDOM}};
  tlbExec_io_in_bits_r_size_p = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  toggle_8690_valid_reg = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  tlbExec_io_in_bits_r_cmd_p = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  toggle_8693_valid_reg = _RAND_32[3:0];
  _RAND_33 = {1{`RANDOM}};
  tlbExec_io_in_bits_r_wmask_p = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  toggle_8697_valid_reg = _RAND_34[7:0];
  _RAND_35 = {2{`RANDOM}};
  tlbExec_io_in_bits_r_wdata_p = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  toggle_8705_valid_reg = _RAND_36[63:0];
  _RAND_37 = {1{`RANDOM}};
  valid_1_p = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  toggle_8769_valid_reg = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  tlbEmpty_io_in_bits_r_addr_p = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  toggle_8770_valid_reg = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  tlbEmpty_io_in_bits_r_size_p = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  toggle_8802_valid_reg = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  tlbEmpty_io_in_bits_r_cmd_p = _RAND_43[3:0];
  _RAND_44 = {1{`RANDOM}};
  toggle_8805_valid_reg = _RAND_44[3:0];
  _RAND_45 = {1{`RANDOM}};
  tlbEmpty_io_in_bits_r_wmask_p = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  toggle_8809_valid_reg = _RAND_46[7:0];
  _RAND_47 = {2{`RANDOM}};
  tlbEmpty_io_in_bits_r_wdata_p = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  toggle_8817_valid_reg = _RAND_48[63:0];
  _RAND_49 = {1{`RANDOM}};
  alreadyOutFinish_p = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  toggle_8881_valid_reg = _RAND_50[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(r_0_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[39]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[40]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[41]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[42]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[43]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[44]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[45]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[46]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[47]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[48]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[49]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[50]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[51]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[52]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[53]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[54]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[55]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[56]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[57]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[58]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[59]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[60]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[61]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[62]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[63]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[64]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[65]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[66]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[67]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[68]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[69]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[70]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[71]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[72]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[73]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[74]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[75]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[76]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[77]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[78]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[79]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[80]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[81]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[82]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[83]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[84]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[85]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[86]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[87]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[88]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[89]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[90]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[91]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[92]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[93]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[94]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[95]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[96]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[97]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[98]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[99]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[100]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[101]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[102]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[103]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[104]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[105]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[106]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[107]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[108]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[109]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[110]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[111]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[112]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[113]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[114]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[115]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[116]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[117]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[118]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[119]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[120]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[121]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[122]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[123]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[124]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[125]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[126]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[127]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[128]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[129]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[130]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[131]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[132]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[133]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[134]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[135]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[136]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[137]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[138]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[139]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[140]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[141]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[142]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[143]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_0_t[144]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[39]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[40]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[41]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[42]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[43]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[44]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[45]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[46]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[47]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[48]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[49]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[50]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[51]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[52]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[53]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[54]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[55]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[56]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[57]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[58]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[59]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[60]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[61]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[62]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[63]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[64]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[65]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[66]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[67]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[68]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[69]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[70]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[71]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[72]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[73]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[74]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[75]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[76]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[77]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[78]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[79]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[80]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[81]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[82]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[83]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[84]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[85]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[86]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[87]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[88]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[89]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[90]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[91]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[92]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[93]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[94]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[95]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[96]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[97]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[98]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[99]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[100]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[101]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[102]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[103]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[104]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[105]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[106]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[107]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[108]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[109]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[110]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[111]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[112]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[113]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[114]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[115]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[116]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[117]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[118]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[119]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[120]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[121]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[122]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[123]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[124]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[125]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[126]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[127]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[128]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[129]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[130]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[131]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[132]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[133]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[134]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[135]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[136]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[137]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[138]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[139]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[140]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[141]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[142]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[143]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_1_t[144]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[39]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[40]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[41]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[42]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[43]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[44]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[45]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[46]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[47]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[48]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[49]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[50]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[51]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[52]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[53]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[54]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[55]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[56]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[57]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[58]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[59]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[60]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[61]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[62]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[63]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[64]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[65]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[66]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[67]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[68]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[69]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[70]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[71]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[72]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[73]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[74]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[75]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[76]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[77]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[78]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[79]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[80]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[81]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[82]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[83]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[84]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[85]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[86]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[87]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[88]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[89]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[90]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[91]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[92]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[93]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[94]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[95]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[96]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[97]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[98]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[99]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[100]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[101]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[102]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[103]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[104]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[105]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[106]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[107]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[108]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[109]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[110]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[111]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[112]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[113]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[114]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[115]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[116]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[117]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[118]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[119]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[120]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[121]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[122]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[123]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[124]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[125]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[126]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[127]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[128]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[129]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[130]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[131]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[132]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[133]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[134]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[135]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[136]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[137]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[138]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[139]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[140]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[141]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[142]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[143]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_2_t[144]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[39]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[40]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[41]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[42]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[43]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[44]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[45]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[46]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[47]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[48]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[49]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[50]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[51]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[52]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[53]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[54]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[55]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[56]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[57]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[58]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[59]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[60]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[61]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[62]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[63]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[64]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[65]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[66]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[67]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[68]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[69]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[70]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[71]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[72]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[73]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[74]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[75]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[76]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[77]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[78]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[79]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[80]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[81]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[82]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[83]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[84]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[85]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[86]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[87]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[88]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[89]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[90]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[91]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[92]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[93]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[94]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[95]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[96]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[97]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[98]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[99]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[100]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[101]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[102]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[103]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[104]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[105]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[106]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[107]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[108]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[109]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[110]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[111]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[112]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[113]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[114]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[115]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[116]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[117]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[118]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[119]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[120]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[121]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[122]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[123]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[124]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[125]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[126]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[127]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[128]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[129]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[130]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[131]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[132]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[133]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[134]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[135]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[136]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[137]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[138]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[139]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[140]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[141]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[142]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[143]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(r_3_t[144]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 96:29]
    end
    //
    if (enToggle_past) begin
      cover(valid_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 107:24]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_addr_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_size_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_size_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_size_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_cmd_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_cmd_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_cmd_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_cmd_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wmask_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wmask_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wmask_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wmask_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wmask_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wmask_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wmask_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wmask_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[0]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[1]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[2]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[3]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[4]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[5]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[6]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[7]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[8]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[9]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[10]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[11]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[12]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[13]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[14]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[15]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[16]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[17]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[18]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[19]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[20]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[21]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[22]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[23]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[24]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[25]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[26]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[27]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[28]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[29]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[30]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[31]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[32]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[33]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[34]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[35]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[36]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[37]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[38]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[39]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[40]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[41]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[42]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[43]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[44]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[45]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[46]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[47]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[48]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[49]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[50]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[51]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[52]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[53]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[54]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[55]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[56]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[57]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[58]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[59]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[60]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[61]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[62]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbExec_io_in_bits_r_wdata_t[63]); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 113:28]
    end
    //
    if (enToggle_past) begin
      cover(valid_1_t); // @[src/main/scala/utils/Pipeline.scala 24:24]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[5]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[6]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[7]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[8]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[9]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[10]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[11]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[12]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[13]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[14]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[15]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[16]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[17]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[18]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[19]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[20]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[21]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[22]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[23]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[24]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[25]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[26]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[27]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[28]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[29]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[30]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_addr_t[31]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_size_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_size_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_size_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_cmd_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_cmd_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_cmd_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_cmd_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wmask_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wmask_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wmask_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wmask_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wmask_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wmask_t[5]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wmask_t[6]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wmask_t[7]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[0]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[1]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[2]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[3]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[4]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[5]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[6]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[7]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[8]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[9]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[10]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[11]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[12]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[13]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[14]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[15]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[16]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[17]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[18]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[19]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[20]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[21]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[22]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[23]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[24]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[25]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[26]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[27]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[28]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[29]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[30]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[31]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[32]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[33]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[34]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[35]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[36]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[37]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[38]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[39]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[40]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[41]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[42]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[43]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[44]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[45]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[46]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[47]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[48]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[49]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[50]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[51]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[52]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[53]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[54]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[55]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[56]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[57]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[58]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[59]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[60]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[61]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[62]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(tlbEmpty_io_in_bits_r_wdata_t[63]); // @[src/main/scala/utils/Pipeline.scala 30:28]
    end
    //
    if (enToggle_past) begin
      cover(alreadyOutFinish_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 176:37]
    end
  end
endmodule
module PTERequestFilter_1(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input         io_out_req_ready, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output        io_out_req_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input         io_out_resp_valid, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input  [63:0] io_out_resp_bits_rdata, // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
  input         io_u // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 549:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
  wire  isLegal = |(io_in_req_bits_addr >= 32'h80000000); // @[src/main/scala/nutcore/NutCore.scala 70:67]
  wire  _hasInflight_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [7:0] _io_in_resp_bits_rdata_T = {3'h7,io_u,4'hf}; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 570:33]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  hasInflight_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
  wire  hasInflight_t = hasInflight ^ hasInflight_p; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
  wire  toggle_8882_clock;
  wire  toggle_8882_reset;
  wire  toggle_8882_valid;
  reg  toggle_8882_valid_reg;
  GEN_w1_toggle #(.COVER_INDEX(8882)) toggle_8882 (
    .clock(toggle_8882_clock),
    .reset(toggle_8882_reset),
    .valid(toggle_8882_valid)
  );
  assign io_in_req_ready = isLegal ? io_out_req_ready : ~hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 562:25]
  assign io_in_resp_valid = ~io_out_resp_valid & hasInflight | io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10 566:44 567:22]
  assign io_in_resp_bits_rdata = ~io_out_resp_valid & hasInflight ? {{56'd0}, _io_in_resp_bits_rdata_T} :
    io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10 566:44 570:27]
  assign io_out_req_valid = io_in_req_valid & isLegal; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 561:39]
  assign io_out_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10]
  assign io_out_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10]
  assign io_out_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 556:10]
  assign toggle_8882_clock = clock;
  assign toggle_8882_reset = reset;
  assign toggle_8882_valid = hasInflight ^ toggle_8882_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
      hasInflight <= 1'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
    end else if (~io_out_resp_valid & hasInflight) begin // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 566:44]
      hasInflight <= 1'h0;
    end else begin
      hasInflight <= _hasInflight_T & ~isLegal; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 564:15]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    hasInflight_p <= hasInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
    toggle_8882_valid_reg <= hasInflight;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  hasInflight = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  hasInflight_p = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  toggle_8882_valid_reg = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(hasInflight_t); // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 559:28]
    end
  end
endmodule
module Cache_fake_1(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_in_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [2:0]  io_in_req_bits_size, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_in_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_out_mem_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_out_mem_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [31:0] io_out_mem_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [2:0]  io_out_mem_req_bits_size, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [3:0]  io_out_mem_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [7:0]  io_out_mem_req_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [63:0] io_out_mem_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_out_mem_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_out_mem_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [3:0]  io_out_mem_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [63:0] io_out_mem_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_mmio_req_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_mmio_req_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [3:0]  io_mmio_req_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [7:0]  io_mmio_req_bits_wmask, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output [63:0] io_mmio_req_bits_wdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        io_mmio_resp_ready, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input         io_mmio_resp_valid, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [3:0]  io_mmio_resp_bits_cmd, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  input  [63:0] io_mmio_resp_bits_rdata, // @[src/main/scala/nutcore/mem/Cache.scala 124:14]
  output        ismmio_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
  wire [31:0] _ismmio_T = io_in_req_bits_addr ^ 32'h30000000; // @[src/main/scala/nutcore/NutCore.scala 114:11]
  wire  _ismmio_T_2 = _ismmio_T[31:28] == 4'h0; // @[src/main/scala/nutcore/NutCore.scala 114:44]
  wire [31:0] _ismmio_T_3 = io_in_req_bits_addr ^ 32'h40000000; // @[src/main/scala/nutcore/NutCore.scala 114:11]
  wire  _ismmio_T_5 = _ismmio_T_3[31:30] == 2'h0; // @[src/main/scala/nutcore/NutCore.scala 114:44]
  wire  ismmio = _ismmio_T_2 | _ismmio_T_5; // @[src/main/scala/nutcore/NutCore.scala 115:15]
  wire  _ismmioRec_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  ismmioRec; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
  reg  alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
  wire  _GEN_3 = io_in_resp_valid | alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 570:{33,33,33}]
  wire  _T_11 = io_out_mem_req_ready & io_out_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_13 = io_out_mem_resp_ready & io_out_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _GEN_6 = _T_13 ? 3'h5 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 581:{37,45}]
  wire  _T_15 = io_mmio_req_ready & io_mmio_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _GEN_7 = _T_15 ? 3'h4 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 584:{33,41}]
  wire  _T_17 = io_mmio_resp_ready & io_mmio_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _GEN_8 = _T_17 | alreadyOutFire ? 3'h5 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 587:{52,60}]
  wire [2:0] _GEN_9 = _GEN_3 ? 3'h0 : state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22 590:{63,71}]
  wire [2:0] _GEN_10 = 3'h5 == state ? _GEN_9 : state; // @[src/main/scala/nutcore/mem/Cache.scala 572:18 558:22]
  wire [2:0] _GEN_11 = 3'h4 == state ? _GEN_8 : _GEN_10; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  wire [2:0] _GEN_12 = 3'h3 == state ? _GEN_7 : _GEN_11; // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
  reg [31:0] reqaddr; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
  reg [3:0] cmd; // @[src/main/scala/nutcore/mem/Cache.scala 595:22]
  reg [2:0] size; // @[src/main/scala/nutcore/mem/Cache.scala 596:23]
  reg [63:0] wdata; // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
  reg [7:0] wmask; // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
  reg [63:0] mmiordata; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
  reg [3:0] mmiocmd; // @[src/main/scala/nutcore/mem/Cache.scala 604:26]
  reg [63:0] memrdata; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
  reg [3:0] memcmd; // @[src/main/scala/nutcore/mem/Cache.scala 606:25]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [2:0] state_p; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
  wire [2:0] state_t = state ^ state_p; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
  wire  toggle_8883_clock;
  wire  toggle_8883_reset;
  wire [2:0] toggle_8883_valid;
  reg [2:0] toggle_8883_valid_reg;
  reg  ismmioRec_p; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
  wire  ismmioRec_t = ismmioRec ^ ismmioRec_p; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
  wire  toggle_8886_clock;
  wire  toggle_8886_reset;
  wire  toggle_8886_valid;
  reg  toggle_8886_valid_reg;
  reg  alreadyOutFire_p; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
  wire  alreadyOutFire_t = alreadyOutFire ^ alreadyOutFire_p; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
  wire  toggle_8887_clock;
  wire  toggle_8887_reset;
  wire  toggle_8887_valid;
  reg  toggle_8887_valid_reg;
  reg [31:0] reqaddr_p; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
  wire [31:0] reqaddr_t = reqaddr ^ reqaddr_p; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
  wire  toggle_8888_clock;
  wire  toggle_8888_reset;
  wire [31:0] toggle_8888_valid;
  reg [31:0] toggle_8888_valid_reg;
  reg [3:0] cmd_p; // @[src/main/scala/nutcore/mem/Cache.scala 595:22]
  wire [3:0] cmd_t = cmd ^ cmd_p; // @[src/main/scala/nutcore/mem/Cache.scala 595:22]
  wire  toggle_8920_clock;
  wire  toggle_8920_reset;
  wire [3:0] toggle_8920_valid;
  reg [3:0] toggle_8920_valid_reg;
  reg [2:0] size_p; // @[src/main/scala/nutcore/mem/Cache.scala 596:23]
  wire [2:0] size_t = size ^ size_p; // @[src/main/scala/nutcore/mem/Cache.scala 596:23]
  wire  toggle_8924_clock;
  wire  toggle_8924_reset;
  wire [2:0] toggle_8924_valid;
  reg [2:0] toggle_8924_valid_reg;
  reg [63:0] wdata_p; // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
  wire [63:0] wdata_t = wdata ^ wdata_p; // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
  wire  toggle_8927_clock;
  wire  toggle_8927_reset;
  wire [63:0] toggle_8927_valid;
  reg [63:0] toggle_8927_valid_reg;
  reg [7:0] wmask_p; // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
  wire [7:0] wmask_t = wmask ^ wmask_p; // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
  wire  toggle_8991_clock;
  wire  toggle_8991_reset;
  wire [7:0] toggle_8991_valid;
  reg [7:0] toggle_8991_valid_reg;
  reg [63:0] mmiordata_p; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
  wire [63:0] mmiordata_t = mmiordata ^ mmiordata_p; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
  wire  toggle_8999_clock;
  wire  toggle_8999_reset;
  wire [63:0] toggle_8999_valid;
  reg [63:0] toggle_8999_valid_reg;
  reg [3:0] mmiocmd_p; // @[src/main/scala/nutcore/mem/Cache.scala 604:26]
  wire [3:0] mmiocmd_t = mmiocmd ^ mmiocmd_p; // @[src/main/scala/nutcore/mem/Cache.scala 604:26]
  wire  toggle_9063_clock;
  wire  toggle_9063_reset;
  wire [3:0] toggle_9063_valid;
  reg [3:0] toggle_9063_valid_reg;
  reg [63:0] memrdata_p; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
  wire [63:0] memrdata_t = memrdata ^ memrdata_p; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
  wire  toggle_9067_clock;
  wire  toggle_9067_reset;
  wire [63:0] toggle_9067_valid;
  reg [63:0] toggle_9067_valid_reg;
  reg [3:0] memcmd_p; // @[src/main/scala/nutcore/mem/Cache.scala 606:25]
  wire [3:0] memcmd_t = memcmd ^ memcmd_p; // @[src/main/scala/nutcore/mem/Cache.scala 606:25]
  wire  toggle_9131_clock;
  wire  toggle_9131_reset;
  wire [3:0] toggle_9131_valid;
  reg [3:0] toggle_9131_valid_reg;
  GEN_w3_toggle #(.COVER_INDEX(8883)) toggle_8883 (
    .clock(toggle_8883_clock),
    .reset(toggle_8883_reset),
    .valid(toggle_8883_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(8886)) toggle_8886 (
    .clock(toggle_8886_clock),
    .reset(toggle_8886_reset),
    .valid(toggle_8886_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(8887)) toggle_8887 (
    .clock(toggle_8887_clock),
    .reset(toggle_8887_reset),
    .valid(toggle_8887_valid)
  );
  GEN_w32_toggle #(.COVER_INDEX(8888)) toggle_8888 (
    .clock(toggle_8888_clock),
    .reset(toggle_8888_reset),
    .valid(toggle_8888_valid)
  );
  GEN_w4_toggle #(.COVER_INDEX(8920)) toggle_8920 (
    .clock(toggle_8920_clock),
    .reset(toggle_8920_reset),
    .valid(toggle_8920_valid)
  );
  GEN_w3_toggle #(.COVER_INDEX(8924)) toggle_8924 (
    .clock(toggle_8924_clock),
    .reset(toggle_8924_reset),
    .valid(toggle_8924_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(8927)) toggle_8927 (
    .clock(toggle_8927_clock),
    .reset(toggle_8927_reset),
    .valid(toggle_8927_valid)
  );
  GEN_w8_toggle #(.COVER_INDEX(8991)) toggle_8991 (
    .clock(toggle_8991_clock),
    .reset(toggle_8991_reset),
    .valid(toggle_8991_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(8999)) toggle_8999 (
    .clock(toggle_8999_clock),
    .reset(toggle_8999_reset),
    .valid(toggle_8999_valid)
  );
  GEN_w4_toggle #(.COVER_INDEX(9063)) toggle_9063 (
    .clock(toggle_9063_clock),
    .reset(toggle_9063_reset),
    .valid(toggle_9063_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(9067)) toggle_9067 (
    .clock(toggle_9067_clock),
    .reset(toggle_9067_reset),
    .valid(toggle_9067_valid)
  );
  GEN_w4_toggle #(.COVER_INDEX(9131)) toggle_9131 (
    .clock(toggle_9131_clock),
    .reset(toggle_9131_reset),
    .valid(toggle_9131_valid)
  );
  assign io_in_req_ready = state == 3'h0; // @[src/main/scala/nutcore/mem/Cache.scala 600:29]
  assign io_in_resp_valid = state == 3'h5; // @[src/main/scala/nutcore/mem/Cache.scala 601:30]
  assign io_in_resp_bits_cmd = ismmioRec ? mmiocmd : memcmd; // @[src/main/scala/nutcore/mem/Cache.scala 609:29]
  assign io_in_resp_bits_rdata = ismmioRec ? mmiordata : memrdata; // @[src/main/scala/nutcore/mem/Cache.scala 608:31]
  assign io_out_mem_req_valid = state == 3'h1; // @[src/main/scala/nutcore/mem/Cache.scala 617:34]
  assign io_out_mem_req_bits_addr = reqaddr; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_out_mem_req_bits_size = size; // @[src/main/scala/bus/simplebus/SimpleBus.scala 66:15]
  assign io_out_mem_req_bits_cmd = cmd; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io_out_mem_req_bits_wmask = wmask; // @[src/main/scala/bus/simplebus/SimpleBus.scala 68:16]
  assign io_out_mem_req_bits_wdata = wdata; // @[src/main/scala/bus/simplebus/SimpleBus.scala 67:16]
  assign io_out_mem_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 618:25]
  assign io_mmio_req_valid = state == 3'h3; // @[src/main/scala/nutcore/mem/Cache.scala 623:31]
  assign io_mmio_req_bits_addr = reqaddr; // @[src/main/scala/bus/simplebus/SimpleBus.scala 64:15]
  assign io_mmio_req_bits_cmd = cmd; // @[src/main/scala/bus/simplebus/SimpleBus.scala 65:14]
  assign io_mmio_req_bits_wmask = wmask; // @[src/main/scala/bus/simplebus/SimpleBus.scala 68:16]
  assign io_mmio_req_bits_wdata = wdata; // @[src/main/scala/bus/simplebus/SimpleBus.scala 67:16]
  assign io_mmio_resp_ready = 1'h1; // @[src/main/scala/nutcore/mem/Cache.scala 624:22]
  assign ismmio_0 = ismmio;
  assign toggle_8883_clock = clock;
  assign toggle_8883_reset = reset;
  assign toggle_8883_valid = state ^ toggle_8883_valid_reg;
  assign toggle_8886_clock = clock;
  assign toggle_8886_reset = reset;
  assign toggle_8886_valid = ismmioRec ^ toggle_8886_valid_reg;
  assign toggle_8887_clock = clock;
  assign toggle_8887_reset = reset;
  assign toggle_8887_valid = alreadyOutFire ^ toggle_8887_valid_reg;
  assign toggle_8888_clock = clock;
  assign toggle_8888_reset = reset;
  assign toggle_8888_valid = reqaddr ^ toggle_8888_valid_reg;
  assign toggle_8920_clock = clock;
  assign toggle_8920_reset = reset;
  assign toggle_8920_valid = cmd ^ toggle_8920_valid_reg;
  assign toggle_8924_clock = clock;
  assign toggle_8924_reset = reset;
  assign toggle_8924_valid = size ^ toggle_8924_valid_reg;
  assign toggle_8927_clock = clock;
  assign toggle_8927_reset = reset;
  assign toggle_8927_valid = wdata ^ toggle_8927_valid_reg;
  assign toggle_8991_clock = clock;
  assign toggle_8991_reset = reset;
  assign toggle_8991_valid = wmask ^ toggle_8991_valid_reg;
  assign toggle_8999_clock = clock;
  assign toggle_8999_reset = reset;
  assign toggle_8999_valid = mmiordata ^ toggle_8999_valid_reg;
  assign toggle_9063_clock = clock;
  assign toggle_9063_reset = reset;
  assign toggle_9063_valid = mmiocmd ^ toggle_9063_valid_reg;
  assign toggle_9067_clock = clock;
  assign toggle_9067_reset = reset;
  assign toggle_9067_valid = memrdata ^ toggle_9067_valid_reg;
  assign toggle_9131_clock = clock;
  assign toggle_9131_reset = reset;
  assign toggle_9131_valid = memcmd ^ toggle_9131_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
      state <= 3'h0; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 575:47]
        if (ismmio) begin // @[src/main/scala/nutcore/mem/Cache.scala 575:61]
          state <= 3'h3;
        end else begin
          state <= 3'h1;
        end
      end
    end else if (3'h1 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      if (_T_11) begin // @[src/main/scala/nutcore/mem/Cache.scala 578:36]
        state <= 3'h2; // @[src/main/scala/nutcore/mem/Cache.scala 578:44]
      end
    end else if (3'h2 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      state <= _GEN_6;
    end else begin
      state <= _GEN_12;
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
      ismmioRec <= ismmio; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
    end
    if (reset) begin // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
    end else if (3'h0 == state) begin // @[src/main/scala/nutcore/mem/Cache.scala 572:18]
      alreadyOutFire <= 1'h0; // @[src/main/scala/nutcore/mem/Cache.scala 574:22]
    end else begin
      alreadyOutFire <= _GEN_3;
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
      reqaddr <= io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 595:22]
      cmd <= io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 595:22]
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 596:23]
      size <= io_in_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 596:23]
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
      wdata <= io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    if (_ismmioRec_T) begin // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
      wmask <= io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
    end
    if (_T_17) begin // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
      mmiordata <= io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    if (_T_17) begin // @[src/main/scala/nutcore/mem/Cache.scala 604:26]
      mmiocmd <= io_mmio_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 604:26]
    end
    if (_T_13) begin // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
      memrdata <= io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    if (_T_13) begin // @[src/main/scala/nutcore/mem/Cache.scala 606:25]
      memcmd <= io_out_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 606:25]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    state_p <= state; // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
    toggle_8883_valid_reg <= state;
    ismmioRec_p <= ismmioRec; // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
    toggle_8886_valid_reg <= ismmioRec;
    alreadyOutFire_p <= alreadyOutFire; // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
    toggle_8887_valid_reg <= alreadyOutFire;
    reqaddr_p <= reqaddr; // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    toggle_8888_valid_reg <= reqaddr;
    cmd_p <= cmd; // @[src/main/scala/nutcore/mem/Cache.scala 595:22]
    toggle_8920_valid_reg <= cmd;
    size_p <= size; // @[src/main/scala/nutcore/mem/Cache.scala 596:23]
    toggle_8924_valid_reg <= size;
    wdata_p <= wdata; // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    toggle_8927_valid_reg <= wdata;
    wmask_p <= wmask; // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
    toggle_8991_valid_reg <= wmask;
    mmiordata_p <= mmiordata; // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    toggle_8999_valid_reg <= mmiordata;
    mmiocmd_p <= mmiocmd; // @[src/main/scala/nutcore/mem/Cache.scala 604:26]
    toggle_9063_valid_reg <= mmiocmd;
    memrdata_p <= memrdata; // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    toggle_9067_valid_reg <= memrdata;
    memcmd_p <= memcmd; // @[src/main/scala/nutcore/mem/Cache.scala 606:25]
    toggle_9131_valid_reg <= memcmd;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  ismmioRec = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  alreadyOutFire = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  reqaddr = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  cmd = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  size = _RAND_5[2:0];
  _RAND_6 = {2{`RANDOM}};
  wdata = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  wmask = _RAND_7[7:0];
  _RAND_8 = {2{`RANDOM}};
  mmiordata = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  mmiocmd = _RAND_9[3:0];
  _RAND_10 = {2{`RANDOM}};
  memrdata = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  memcmd = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  state_p = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  toggle_8883_valid_reg = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  ismmioRec_p = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  toggle_8886_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  alreadyOutFire_p = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  toggle_8887_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  reqaddr_p = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  toggle_8888_valid_reg = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  cmd_p = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  toggle_8920_valid_reg = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  size_p = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  toggle_8924_valid_reg = _RAND_23[2:0];
  _RAND_24 = {2{`RANDOM}};
  wdata_p = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  toggle_8927_valid_reg = _RAND_25[63:0];
  _RAND_26 = {1{`RANDOM}};
  wmask_p = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  toggle_8991_valid_reg = _RAND_27[7:0];
  _RAND_28 = {2{`RANDOM}};
  mmiordata_p = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  toggle_8999_valid_reg = _RAND_29[63:0];
  _RAND_30 = {1{`RANDOM}};
  mmiocmd_p = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
  toggle_9063_valid_reg = _RAND_31[3:0];
  _RAND_32 = {2{`RANDOM}};
  memrdata_p = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  toggle_9067_valid_reg = _RAND_33[63:0];
  _RAND_34 = {1{`RANDOM}};
  memcmd_p = _RAND_34[3:0];
  _RAND_35 = {1{`RANDOM}};
  toggle_9131_valid_reg = _RAND_35[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(state_t[0]); // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[1]); // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[2]); // @[src/main/scala/nutcore/mem/Cache.scala 558:22]
    end
    //
    if (enToggle_past) begin
      cover(ismmioRec_t); // @[src/main/scala/nutcore/mem/Cache.scala 561:28]
    end
    //
    if (enToggle_past) begin
      cover(alreadyOutFire_t); // @[src/main/scala/nutcore/mem/Cache.scala 570:33]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[0]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[1]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[2]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[3]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[4]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[5]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[6]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[7]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[8]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[9]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[10]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[11]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[12]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[13]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[14]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[15]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[16]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[17]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[18]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[19]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[20]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[21]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[22]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[23]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[24]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[25]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[26]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[27]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[28]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[29]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[30]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(reqaddr_t[31]); // @[src/main/scala/nutcore/mem/Cache.scala 594:26]
    end
    //
    if (enToggle_past) begin
      cover(cmd_t[0]); // @[src/main/scala/nutcore/mem/Cache.scala 595:22]
    end
    //
    if (enToggle_past) begin
      cover(cmd_t[1]); // @[src/main/scala/nutcore/mem/Cache.scala 595:22]
    end
    //
    if (enToggle_past) begin
      cover(cmd_t[2]); // @[src/main/scala/nutcore/mem/Cache.scala 595:22]
    end
    //
    if (enToggle_past) begin
      cover(cmd_t[3]); // @[src/main/scala/nutcore/mem/Cache.scala 595:22]
    end
    //
    if (enToggle_past) begin
      cover(size_t[0]); // @[src/main/scala/nutcore/mem/Cache.scala 596:23]
    end
    //
    if (enToggle_past) begin
      cover(size_t[1]); // @[src/main/scala/nutcore/mem/Cache.scala 596:23]
    end
    //
    if (enToggle_past) begin
      cover(size_t[2]); // @[src/main/scala/nutcore/mem/Cache.scala 596:23]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[0]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[1]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[2]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[3]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[4]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[5]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[6]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[7]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[8]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[9]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[10]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[11]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[12]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[13]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[14]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[15]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[16]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[17]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[18]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[19]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[20]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[21]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[22]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[23]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[24]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[25]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[26]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[27]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[28]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[29]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[30]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[31]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[32]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[33]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[34]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[35]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[36]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[37]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[38]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[39]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[40]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[41]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[42]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[43]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[44]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[45]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[46]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[47]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[48]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[49]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[50]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[51]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[52]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[53]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[54]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[55]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[56]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[57]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[58]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[59]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[60]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[61]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[62]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wdata_t[63]); // @[src/main/scala/nutcore/mem/Cache.scala 597:24]
    end
    //
    if (enToggle_past) begin
      cover(wmask_t[0]); // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
    end
    //
    if (enToggle_past) begin
      cover(wmask_t[1]); // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
    end
    //
    if (enToggle_past) begin
      cover(wmask_t[2]); // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
    end
    //
    if (enToggle_past) begin
      cover(wmask_t[3]); // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
    end
    //
    if (enToggle_past) begin
      cover(wmask_t[4]); // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
    end
    //
    if (enToggle_past) begin
      cover(wmask_t[5]); // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
    end
    //
    if (enToggle_past) begin
      cover(wmask_t[6]); // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
    end
    //
    if (enToggle_past) begin
      cover(wmask_t[7]); // @[src/main/scala/nutcore/mem/Cache.scala 598:24]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[0]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[1]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[2]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[3]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[4]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[5]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[6]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[7]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[8]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[9]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[10]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[11]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[12]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[13]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[14]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[15]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[16]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[17]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[18]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[19]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[20]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[21]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[22]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[23]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[24]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[25]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[26]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[27]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[28]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[29]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[30]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[31]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[32]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[33]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[34]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[35]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[36]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[37]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[38]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[39]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[40]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[41]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[42]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[43]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[44]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[45]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[46]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[47]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[48]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[49]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[50]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[51]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[52]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[53]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[54]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[55]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[56]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[57]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[58]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[59]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[60]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[61]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[62]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiordata_t[63]); // @[src/main/scala/nutcore/mem/Cache.scala 603:28]
    end
    //
    if (enToggle_past) begin
      cover(mmiocmd_t[0]); // @[src/main/scala/nutcore/mem/Cache.scala 604:26]
    end
    //
    if (enToggle_past) begin
      cover(mmiocmd_t[1]); // @[src/main/scala/nutcore/mem/Cache.scala 604:26]
    end
    //
    if (enToggle_past) begin
      cover(mmiocmd_t[2]); // @[src/main/scala/nutcore/mem/Cache.scala 604:26]
    end
    //
    if (enToggle_past) begin
      cover(mmiocmd_t[3]); // @[src/main/scala/nutcore/mem/Cache.scala 604:26]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[0]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[1]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[2]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[3]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[4]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[5]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[6]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[7]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[8]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[9]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[10]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[11]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[12]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[13]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[14]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[15]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[16]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[17]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[18]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[19]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[20]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[21]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[22]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[23]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[24]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[25]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[26]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[27]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[28]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[29]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[30]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[31]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[32]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[33]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[34]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[35]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[36]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[37]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[38]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[39]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[40]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[41]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[42]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[43]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[44]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[45]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[46]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[47]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[48]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[49]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[50]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[51]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[52]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[53]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[54]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[55]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[56]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[57]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[58]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[59]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[60]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[61]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[62]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memrdata_t[63]); // @[src/main/scala/nutcore/mem/Cache.scala 605:27]
    end
    //
    if (enToggle_past) begin
      cover(memcmd_t[0]); // @[src/main/scala/nutcore/mem/Cache.scala 606:25]
    end
    //
    if (enToggle_past) begin
      cover(memcmd_t[1]); // @[src/main/scala/nutcore/mem/Cache.scala 606:25]
    end
    //
    if (enToggle_past) begin
      cover(memcmd_t[2]); // @[src/main/scala/nutcore/mem/Cache.scala 606:25]
    end
    //
    if (enToggle_past) begin
      cover(memcmd_t[3]); // @[src/main/scala/nutcore/mem/Cache.scala 606:25]
    end
  end
endmodule
module NutCore(
  input         clock,
  input         reset,
  input         io_imem_mem_req_ready, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output        io_imem_mem_req_valid, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [31:0] io_imem_mem_req_bits_addr, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input         io_imem_mem_resp_valid, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input  [63:0] io_imem_mem_resp_bits_rdata, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input         io_dmem_mem_req_ready, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output        io_dmem_mem_req_valid, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [31:0] io_dmem_mem_req_bits_addr, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [2:0]  io_dmem_mem_req_bits_size, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [3:0]  io_dmem_mem_req_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [7:0]  io_dmem_mem_req_bits_wmask, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [63:0] io_dmem_mem_req_bits_wdata, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input         io_dmem_mem_resp_valid, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input  [3:0]  io_dmem_mem_resp_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input  [63:0] io_dmem_mem_resp_bits_rdata, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input         io_mmio_req_ready, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output        io_mmio_req_valid, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [3:0]  io_mmio_req_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [7:0]  io_mmio_req_bits_wmask, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  output [63:0] io_mmio_req_bits_wdata, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input         io_mmio_resp_valid, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input  [3:0]  io_mmio_resp_bits_cmd, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input  [63:0] io_mmio_resp_bits_rdata, // @[src/main/scala/nutcore/NutCore.scala 125:14]
  input         io_extra_meip_0,
  output        isWFI,
  input         io_extra_mtip,
  input         io_extra_msip
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [63:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [63:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [63:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [63:0] _RAND_240;
  reg [63:0] _RAND_241;
  reg [63:0] _RAND_242;
  reg [63:0] _RAND_243;
  reg [63:0] _RAND_244;
  reg [63:0] _RAND_245;
  reg [63:0] _RAND_246;
  reg [63:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [63:0] _RAND_288;
  reg [63:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
`endif // RANDOMIZE_REG_INIT
  wire  frontend_clock; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_reset; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_imem_req_ready; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_imem_req_valid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [38:0] frontend_io_imem_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [86:0] frontend_io_imem_req_bits_user; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_imem_resp_ready; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_imem_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [63:0] frontend_io_imem_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [86:0] frontend_io_imem_resp_bits_user; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_ready; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_valid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [63:0] frontend_io_out_0_bits_cf_instr; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [38:0] frontend_io_out_0_bits_cf_pc; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [38:0] frontend_io_out_0_bits_cf_pnpc; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [3:0] frontend_io_out_0_bits_cf_brIdx; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [2:0] frontend_io_out_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [6:0] frontend_io_out_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_out_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [63:0] frontend_io_out_0_bits_data_imm; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [3:0] frontend_io_flushVec; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [38:0] frontend_io_redirect_target; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_redirect_valid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_iaf; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_sfence_vma_invalid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_io_wfi_invalid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_REG_valid; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [38:0] frontend_REG_pc; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_REG_isMissPredict; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [38:0] frontend_REG_actualTarget; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [6:0] frontend_REG_fuOpType; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [1:0] frontend_REG_btbType; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_REG_isRVC; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_isWFI; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_flushICache; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  frontend_flushTLB; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire [11:0] frontend_intrVecIDU; // @[src/main/scala/nutcore/NutCore.scala 131:34]
  wire  backend_clock; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_reset; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_ready; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_valid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [63:0] backend_io_in_0_bits_cf_instr; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [38:0] backend_io_in_0_bits_cf_pc; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [38:0] backend_io_in_0_bits_cf_pnpc; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_exceptionVec_1; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_exceptionVec_2; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_exceptionVec_12; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_intrVec_1; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_intrVec_3; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_intrVec_5; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_intrVec_7; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_intrVec_9; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_intrVec_11; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [3:0] backend_io_in_0_bits_cf_brIdx; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_cf_crossBoundaryFault; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_ctrl_src1Type; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_ctrl_src2Type; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [2:0] backend_io_in_0_bits_ctrl_fuType; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [6:0] backend_io_in_0_bits_ctrl_fuOpType; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [4:0] backend_io_in_0_bits_ctrl_rfSrc1; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [4:0] backend_io_in_0_bits_ctrl_rfSrc2; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_ctrl_rfWen; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [4:0] backend_io_in_0_bits_ctrl_rfDest; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_in_0_bits_ctrl_isNutCoreTrap; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [63:0] backend_io_in_0_bits_data_imm; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [1:0] backend_io_flush; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_dmem_req_ready; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_dmem_req_valid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [38:0] backend_io_dmem_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [2:0] backend_io_dmem_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [3:0] backend_io_dmem_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [7:0] backend_io_dmem_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [63:0] backend_io_dmem_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_dmem_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [63:0] backend_io_dmem_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [1:0] backend_io_memMMU_imem_priviledgeMode; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [1:0] backend_io_memMMU_dmem_priviledgeMode; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_memMMU_dmem_status_sum; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_memMMU_dmem_status_mxr; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_memMMU_dmem_loadPF; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_memMMU_dmem_storePF; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_memMMU_dmem_laf; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_memMMU_dmem_saf; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_sfence_vma_invalid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_wfi_invalid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [38:0] backend_io_redirect_target; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_redirect_valid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_lr; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_extra_meip_0; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_scInflight; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_REG_valid; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [38:0] backend_REG_pc; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_REG_isMissPredict; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [38:0] backend_REG_actualTarget; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [6:0] backend_REG_fuOpType; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [1:0] backend_REG_btbType; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_REG_isRVC; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_amoReq; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [63:0] backend_lrAddr; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [55:0] backend_paddr; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [63:0] backend_satp; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend__T_12; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_scIsSuccess; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_extra_mtip; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_flushICache; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_vmEnable; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_flushTLB; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire [11:0] backend_intrVecIDU; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_tlbFinish; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_ismmio; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend__T_13_0; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  backend_io_extra_msip; // @[src/main/scala/nutcore/NutCore.scala 174:25]
  wire  mmioXbar_clock; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_reset; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_in_0_req_ready; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_in_0_req_valid; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [31:0] mmioXbar_io_in_0_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_in_0_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [63:0] mmioXbar_io_in_0_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_in_1_req_ready; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_in_1_req_valid; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [31:0] mmioXbar_io_in_1_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [3:0] mmioXbar_io_in_1_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [7:0] mmioXbar_io_in_1_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [63:0] mmioXbar_io_in_1_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_in_1_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [3:0] mmioXbar_io_in_1_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [63:0] mmioXbar_io_in_1_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_out_req_ready; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_out_req_valid; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [31:0] mmioXbar_io_out_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [3:0] mmioXbar_io_out_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [7:0] mmioXbar_io_out_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [63:0] mmioXbar_io_out_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_out_resp_ready; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  mmioXbar_io_out_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [3:0] mmioXbar_io_out_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire [63:0] mmioXbar_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 178:26]
  wire  dmemXbar_clock; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_reset; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_0_req_ready; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_0_req_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [31:0] dmemXbar_io_in_0_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [2:0] dmemXbar_io_in_0_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [3:0] dmemXbar_io_in_0_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [7:0] dmemXbar_io_in_0_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_in_0_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_0_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_in_0_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_1_req_ready; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_1_req_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [31:0] dmemXbar_io_in_1_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [3:0] dmemXbar_io_in_1_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_in_1_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_1_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_in_1_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_2_req_ready; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_2_req_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [31:0] dmemXbar_io_in_2_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [3:0] dmemXbar_io_in_2_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_in_2_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_in_2_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_in_2_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_out_req_ready; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_out_req_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [31:0] dmemXbar_io_out_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [2:0] dmemXbar_io_out_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [3:0] dmemXbar_io_out_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [7:0] dmemXbar_io_out_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_out_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_out_resp_ready; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  dmemXbar_io_out_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [3:0] dmemXbar_io_out_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire [63:0] dmemXbar_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 179:26]
  wire  itlb_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_in_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [38:0] itlb_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [86:0] itlb_io_in_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_in_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] itlb_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [86:0] itlb_io_in_resp_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [31:0] itlb_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [86:0] itlb_io_out_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_out_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] itlb_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [86:0] itlb_io_out_resp_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [31:0] itlb_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [3:0] itlb_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] itlb_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] itlb_io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_flush; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [1:0] itlb_io_csrMMU_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_io_iaf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] itlb_CSRSATP; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  itlb_MOUFlushTLB; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  filter_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_in_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [31:0] filter_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [3:0] filter_io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [31:0] filter_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [3:0] filter_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_io_u; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  io_imem_cache_clock; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_reset; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_in_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_imem_cache_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [86:0] io_imem_cache_io_in_req_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_in_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_imem_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [86:0] io_imem_cache_io_in_resp_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [1:0] io_imem_cache_io_flush; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_out_mem_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_imem_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_out_mem_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_out_mem_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_imem_cache_io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_mmio_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_imem_cache_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_mmio_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_imem_cache_io_mmio_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_imem_cache_io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  dtlb_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_in_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [38:0] dtlb_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [2:0] dtlb_io_in_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [3:0] dtlb_io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [7:0] dtlb_io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [31:0] dtlb_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [2:0] dtlb_io_out_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [3:0] dtlb_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [7:0] dtlb_io_out_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_mem_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [31:0] dtlb_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [3:0] dtlb_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_mem_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_io_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [1:0] dtlb_io_csrMMU_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_csrMMU_status_sum; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_csrMMU_status_mxr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_csrMMU_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_csrMMU_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_csrMMU_laf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_io_csrMMU_saf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_lr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_scInflight; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_amoReq; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_lrAddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [55:0] dtlb_paddr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire [63:0] dtlb_CSRSATP; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb__T_12_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_scIsSuccess_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_vmEnable_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_MOUFlushTLB; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb_tlbFinish_0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  dtlb__T_13_1; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
  wire  filter_1_clock; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_reset; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_in_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [31:0] filter_1_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [3:0] filter_1_io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_1_io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_1_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_out_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [31:0] filter_1_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [3:0] filter_1_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_1_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_out_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire [63:0] filter_1_io_out_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  filter_1_io_u; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
  wire  io_dmem_cache_clock; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_reset; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_in_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_dmem_cache_io_in_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [2:0] io_dmem_cache_io_in_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_in_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [7:0] io_dmem_cache_io_in_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_in_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_in_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_out_mem_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_dmem_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [2:0] io_dmem_cache_io_out_mem_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_out_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [7:0] io_dmem_cache_io_out_mem_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_out_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_out_mem_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_out_mem_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_out_mem_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_out_mem_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_mmio_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [31:0] io_dmem_cache_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_mmio_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [7:0] io_dmem_cache_io_mmio_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_mmio_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_mmio_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_io_mmio_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [3:0] io_dmem_cache_io_mmio_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire [63:0] io_dmem_cache_io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  wire  io_dmem_cache_ismmio_0; // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
  reg [63:0] dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [3:0] dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [2:0] dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [6:0] dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_0_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_1_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_1_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_1_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [3:0] dataBuffer_1_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [2:0] dataBuffer_1_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [6:0] dataBuffer_1_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_1_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_1_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_1_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_1_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_1_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_2_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_2_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_2_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [3:0] dataBuffer_2_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [2:0] dataBuffer_2_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [6:0] dataBuffer_2_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_2_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_2_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_2_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_2_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_2_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_3_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_3_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [38:0] dataBuffer_3_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [3:0] dataBuffer_3_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [2:0] dataBuffer_3_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [6:0] dataBuffer_3_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_3_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_3_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [4:0] dataBuffer_3_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg  dataBuffer_3_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [63:0] dataBuffer_3_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  reg [1:0] ringBufferHead; // @[src/main/scala/utils/PipelineVector.scala 30:33]
  reg [1:0] ringBufferTail; // @[src/main/scala/utils/PipelineVector.scala 31:33]
  wire [1:0] _ringBufferAllowin_T_1 = ringBufferHead + 2'h1; // @[src/main/scala/utils/PipelineVector.scala 33:63]
  wire [1:0] _ringBufferAllowin_T_4 = ringBufferHead + 2'h2; // @[src/main/scala/utils/PipelineVector.scala 33:63]
  wire  ringBufferAllowin = _ringBufferAllowin_T_1 != ringBufferTail & _ringBufferAllowin_T_4 != ringBufferTail; // @[src/main/scala/utils/PipelineVector.scala 33:124]
  wire  needEnqueue_0 = frontend_io_out_0_valid; // @[src/main/scala/utils/PipelineVector.scala 36:27 37:20]
  wire [1:0] enqueueSize = {{1'd0}, needEnqueue_0}; // @[src/main/scala/utils/PipelineVector.scala 40:44]
  wire  enqueueFire_0 = enqueueSize >= 2'h1; // @[src/main/scala/utils/PipelineVector.scala 41:53]
  wire  enqueueFire_1 = enqueueSize >= 2'h2; // @[src/main/scala/utils/PipelineVector.scala 41:53]
  wire  wen = frontend_io_out_0_ready & frontend_io_out_0_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _T_1 = {{1'd0}, ringBufferHead}; // @[src/main/scala/utils/PipelineVector.scala 45:45]
  wire [63:0] _dataBuffer_T_cf_instr = needEnqueue_0 ? frontend_io_out_0_bits_cf_instr : 64'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [38:0] _dataBuffer_T_cf_pc = needEnqueue_0 ? frontend_io_out_0_bits_cf_pc : 39'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [38:0] _dataBuffer_T_cf_pnpc = needEnqueue_0 ? frontend_io_out_0_bits_cf_pnpc : 39'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [3:0] _dataBuffer_T_cf_brIdx = needEnqueue_0 ? frontend_io_out_0_bits_cf_brIdx : 4'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [2:0] _dataBuffer_T_ctrl_fuType = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_fuType : 3'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [6:0] _dataBuffer_T_ctrl_fuOpType = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_fuOpType : 7'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [4:0] _dataBuffer_T_ctrl_rfSrc1 = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_rfSrc1 : 5'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [4:0] _dataBuffer_T_ctrl_rfSrc2 = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_rfSrc2 : 5'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [4:0] _dataBuffer_T_ctrl_rfDest = needEnqueue_0 ? frontend_io_out_0_bits_ctrl_rfDest : 5'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [63:0] _dataBuffer_T_data_imm = needEnqueue_0 ? frontend_io_out_0_bits_data_imm : 64'h0; // @[src/main/scala/utils/PipelineVector.scala 45:69]
  wire [63:0] _GEN_0 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_instr : dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_1 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_instr : dataBuffer_1_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_2 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_instr : dataBuffer_2_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_3 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_instr : dataBuffer_3_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_4 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_pc : dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_5 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_pc : dataBuffer_1_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_6 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_pc : dataBuffer_2_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_7 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_pc : dataBuffer_3_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_8 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_pnpc : dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_9 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_pnpc : dataBuffer_1_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_10 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_pnpc : dataBuffer_2_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [38:0] _GEN_11 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_pnpc : dataBuffer_3_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_28 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_1 :
    dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_29 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_1 :
    dataBuffer_1_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_30 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_1 :
    dataBuffer_2_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_31 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_1 :
    dataBuffer_3_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_32 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_2 :
    dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_33 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_2 :
    dataBuffer_1_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_34 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_2 :
    dataBuffer_2_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_35 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_2 :
    dataBuffer_3_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_72 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    dataBuffer_0_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_73 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    dataBuffer_1_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_74 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    dataBuffer_2_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_75 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_exceptionVec_12 :
    dataBuffer_3_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_92 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_1 : dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_93 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_1 : dataBuffer_1_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_94 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_1 : dataBuffer_2_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_95 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_1 : dataBuffer_3_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_100 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_3 : dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_101 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_3 : dataBuffer_1_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_102 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_3 : dataBuffer_2_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_103 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_3 : dataBuffer_3_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_108 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_5 : dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_109 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_5 : dataBuffer_1_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_110 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_5 : dataBuffer_2_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_111 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_5 : dataBuffer_3_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_116 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_7 : dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_117 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_7 : dataBuffer_1_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_118 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_7 : dataBuffer_2_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_119 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_7 : dataBuffer_3_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_124 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_9 : dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_125 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_9 : dataBuffer_1_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_126 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_9 : dataBuffer_2_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_127 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_9 : dataBuffer_3_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_132 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_11 : dataBuffer_0_cf_intrVec_11
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_133 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_11 : dataBuffer_1_cf_intrVec_11
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_134 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_11 : dataBuffer_2_cf_intrVec_11
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_135 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_intrVec_11 : dataBuffer_3_cf_intrVec_11
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_136 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_cf_brIdx : dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_137 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_cf_brIdx : dataBuffer_1_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_138 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_cf_brIdx : dataBuffer_2_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [3:0] _GEN_139 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_cf_brIdx : dataBuffer_3_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_144 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_crossBoundaryFault :
    dataBuffer_0_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_145 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_crossBoundaryFault :
    dataBuffer_1_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_146 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_crossBoundaryFault :
    dataBuffer_2_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_147 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_cf_crossBoundaryFault :
    dataBuffer_3_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_160 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src1Type : dataBuffer_0_ctrl_src1Type
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_161 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src1Type : dataBuffer_1_ctrl_src1Type
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_162 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src1Type : dataBuffer_2_ctrl_src1Type
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_163 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src1Type : dataBuffer_3_ctrl_src1Type
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_164 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src2Type : dataBuffer_0_ctrl_src2Type
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_165 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src2Type : dataBuffer_1_ctrl_src2Type
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_166 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src2Type : dataBuffer_2_ctrl_src2Type
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_167 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_src2Type : dataBuffer_3_ctrl_src2Type
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_168 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuType : dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_169 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuType : dataBuffer_1_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_170 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuType : dataBuffer_2_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [2:0] _GEN_171 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuType : dataBuffer_3_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_172 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuOpType : dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_173 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuOpType : dataBuffer_1_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_174 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuOpType : dataBuffer_2_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [6:0] _GEN_175 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_fuOpType : dataBuffer_3_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_176 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc1 : dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_177 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc1 : dataBuffer_1_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_178 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc1 : dataBuffer_2_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_179 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc1 : dataBuffer_3_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_180 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc2 : dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_181 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc2 : dataBuffer_1_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_182 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc2 : dataBuffer_2_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_183 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfSrc2 : dataBuffer_3_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_184 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_rfWen : dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_185 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_rfWen : dataBuffer_1_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_186 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_rfWen : dataBuffer_2_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_187 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_rfWen : dataBuffer_3_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_188 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfDest : dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_189 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfDest : dataBuffer_1_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_190 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfDest : dataBuffer_2_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [4:0] _GEN_191 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_ctrl_rfDest : dataBuffer_3_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_192 = 2'h0 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_isNutCoreTrap :
    dataBuffer_0_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_193 = 2'h1 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_isNutCoreTrap :
    dataBuffer_1_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_194 = 2'h2 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_isNutCoreTrap :
    dataBuffer_2_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire  _GEN_195 = 2'h3 == _T_1[1:0] ? needEnqueue_0 & frontend_io_out_0_bits_ctrl_isNutCoreTrap :
    dataBuffer_3_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_220 = 2'h0 == _T_1[1:0] ? _dataBuffer_T_data_imm : dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_221 = 2'h1 == _T_1[1:0] ? _dataBuffer_T_data_imm : dataBuffer_1_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_222 = 2'h2 == _T_1[1:0] ? _dataBuffer_T_data_imm : dataBuffer_2_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_223 = 2'h3 == _T_1[1:0] ? _dataBuffer_T_data_imm : dataBuffer_3_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:{63,63}]
  wire [63:0] _GEN_224 = enqueueFire_0 ? _GEN_0 : dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_225 = enqueueFire_0 ? _GEN_1 : dataBuffer_1_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_226 = enqueueFire_0 ? _GEN_2 : dataBuffer_2_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_227 = enqueueFire_0 ? _GEN_3 : dataBuffer_3_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_228 = enqueueFire_0 ? _GEN_4 : dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_229 = enqueueFire_0 ? _GEN_5 : dataBuffer_1_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_230 = enqueueFire_0 ? _GEN_6 : dataBuffer_2_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_231 = enqueueFire_0 ? _GEN_7 : dataBuffer_3_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_232 = enqueueFire_0 ? _GEN_8 : dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_233 = enqueueFire_0 ? _GEN_9 : dataBuffer_1_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_234 = enqueueFire_0 ? _GEN_10 : dataBuffer_2_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [38:0] _GEN_235 = enqueueFire_0 ? _GEN_11 : dataBuffer_3_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_252 = enqueueFire_0 ? _GEN_28 : dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_253 = enqueueFire_0 ? _GEN_29 : dataBuffer_1_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_254 = enqueueFire_0 ? _GEN_30 : dataBuffer_2_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_255 = enqueueFire_0 ? _GEN_31 : dataBuffer_3_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_256 = enqueueFire_0 ? _GEN_32 : dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_257 = enqueueFire_0 ? _GEN_33 : dataBuffer_1_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_258 = enqueueFire_0 ? _GEN_34 : dataBuffer_2_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_259 = enqueueFire_0 ? _GEN_35 : dataBuffer_3_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_296 = enqueueFire_0 ? _GEN_72 : dataBuffer_0_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_297 = enqueueFire_0 ? _GEN_73 : dataBuffer_1_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_298 = enqueueFire_0 ? _GEN_74 : dataBuffer_2_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_299 = enqueueFire_0 ? _GEN_75 : dataBuffer_3_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_316 = enqueueFire_0 ? _GEN_92 : dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_317 = enqueueFire_0 ? _GEN_93 : dataBuffer_1_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_318 = enqueueFire_0 ? _GEN_94 : dataBuffer_2_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_319 = enqueueFire_0 ? _GEN_95 : dataBuffer_3_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_324 = enqueueFire_0 ? _GEN_100 : dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_325 = enqueueFire_0 ? _GEN_101 : dataBuffer_1_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_326 = enqueueFire_0 ? _GEN_102 : dataBuffer_2_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_327 = enqueueFire_0 ? _GEN_103 : dataBuffer_3_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_332 = enqueueFire_0 ? _GEN_108 : dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_333 = enqueueFire_0 ? _GEN_109 : dataBuffer_1_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_334 = enqueueFire_0 ? _GEN_110 : dataBuffer_2_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_335 = enqueueFire_0 ? _GEN_111 : dataBuffer_3_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_340 = enqueueFire_0 ? _GEN_116 : dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_341 = enqueueFire_0 ? _GEN_117 : dataBuffer_1_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_342 = enqueueFire_0 ? _GEN_118 : dataBuffer_2_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_343 = enqueueFire_0 ? _GEN_119 : dataBuffer_3_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_348 = enqueueFire_0 ? _GEN_124 : dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_349 = enqueueFire_0 ? _GEN_125 : dataBuffer_1_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_350 = enqueueFire_0 ? _GEN_126 : dataBuffer_2_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_351 = enqueueFire_0 ? _GEN_127 : dataBuffer_3_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_356 = enqueueFire_0 ? _GEN_132 : dataBuffer_0_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_357 = enqueueFire_0 ? _GEN_133 : dataBuffer_1_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_358 = enqueueFire_0 ? _GEN_134 : dataBuffer_2_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_359 = enqueueFire_0 ? _GEN_135 : dataBuffer_3_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_360 = enqueueFire_0 ? _GEN_136 : dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_361 = enqueueFire_0 ? _GEN_137 : dataBuffer_1_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_362 = enqueueFire_0 ? _GEN_138 : dataBuffer_2_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [3:0] _GEN_363 = enqueueFire_0 ? _GEN_139 : dataBuffer_3_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_368 = enqueueFire_0 ? _GEN_144 : dataBuffer_0_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_369 = enqueueFire_0 ? _GEN_145 : dataBuffer_1_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_370 = enqueueFire_0 ? _GEN_146 : dataBuffer_2_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_371 = enqueueFire_0 ? _GEN_147 : dataBuffer_3_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_384 = enqueueFire_0 ? _GEN_160 : dataBuffer_0_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_385 = enqueueFire_0 ? _GEN_161 : dataBuffer_1_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_386 = enqueueFire_0 ? _GEN_162 : dataBuffer_2_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_387 = enqueueFire_0 ? _GEN_163 : dataBuffer_3_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_388 = enqueueFire_0 ? _GEN_164 : dataBuffer_0_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_389 = enqueueFire_0 ? _GEN_165 : dataBuffer_1_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_390 = enqueueFire_0 ? _GEN_166 : dataBuffer_2_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_391 = enqueueFire_0 ? _GEN_167 : dataBuffer_3_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_392 = enqueueFire_0 ? _GEN_168 : dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_393 = enqueueFire_0 ? _GEN_169 : dataBuffer_1_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_394 = enqueueFire_0 ? _GEN_170 : dataBuffer_2_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [2:0] _GEN_395 = enqueueFire_0 ? _GEN_171 : dataBuffer_3_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_396 = enqueueFire_0 ? _GEN_172 : dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_397 = enqueueFire_0 ? _GEN_173 : dataBuffer_1_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_398 = enqueueFire_0 ? _GEN_174 : dataBuffer_2_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [6:0] _GEN_399 = enqueueFire_0 ? _GEN_175 : dataBuffer_3_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_400 = enqueueFire_0 ? _GEN_176 : dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_401 = enqueueFire_0 ? _GEN_177 : dataBuffer_1_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_402 = enqueueFire_0 ? _GEN_178 : dataBuffer_2_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_403 = enqueueFire_0 ? _GEN_179 : dataBuffer_3_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_404 = enqueueFire_0 ? _GEN_180 : dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_405 = enqueueFire_0 ? _GEN_181 : dataBuffer_1_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_406 = enqueueFire_0 ? _GEN_182 : dataBuffer_2_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_407 = enqueueFire_0 ? _GEN_183 : dataBuffer_3_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_408 = enqueueFire_0 ? _GEN_184 : dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_409 = enqueueFire_0 ? _GEN_185 : dataBuffer_1_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_410 = enqueueFire_0 ? _GEN_186 : dataBuffer_2_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_411 = enqueueFire_0 ? _GEN_187 : dataBuffer_3_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_412 = enqueueFire_0 ? _GEN_188 : dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_413 = enqueueFire_0 ? _GEN_189 : dataBuffer_1_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_414 = enqueueFire_0 ? _GEN_190 : dataBuffer_2_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [4:0] _GEN_415 = enqueueFire_0 ? _GEN_191 : dataBuffer_3_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_416 = enqueueFire_0 ? _GEN_192 : dataBuffer_0_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_417 = enqueueFire_0 ? _GEN_193 : dataBuffer_1_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_418 = enqueueFire_0 ? _GEN_194 : dataBuffer_2_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire  _GEN_419 = enqueueFire_0 ? _GEN_195 : dataBuffer_3_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_444 = enqueueFire_0 ? _GEN_220 : dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_445 = enqueueFire_0 ? _GEN_221 : dataBuffer_1_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_446 = enqueueFire_0 ? _GEN_222 : dataBuffer_2_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [63:0] _GEN_447 = enqueueFire_0 ? _GEN_223 : dataBuffer_3_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29 45:29]
  wire [1:0] _T_4 = 2'h1 + ringBufferHead; // @[src/main/scala/utils/PipelineVector.scala 46:45]
  wire [1:0] _ringBufferHead_T_1 = ringBufferHead + enqueueSize; // @[src/main/scala/utils/PipelineVector.scala 47:42]
  wire [63:0] _GEN_1122 = 2'h1 == ringBufferTail ? dataBuffer_1_data_imm : dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_1123 = 2'h2 == ringBufferTail ? dataBuffer_2_data_imm : _GEN_1122; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1150 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_isNutCoreTrap : dataBuffer_0_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1151 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_isNutCoreTrap : _GEN_1150; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1154 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_rfDest : dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1155 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_rfDest : _GEN_1154; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1158 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_rfWen : dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1159 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_rfWen : _GEN_1158; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1162 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_rfSrc2 : dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1163 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_rfSrc2 : _GEN_1162; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1166 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_rfSrc1 : dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [4:0] _GEN_1167 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_rfSrc1 : _GEN_1166; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [6:0] _GEN_1170 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_fuOpType : dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [6:0] _GEN_1171 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_fuOpType : _GEN_1170; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [2:0] _GEN_1174 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_fuType : dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [2:0] _GEN_1175 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_fuType : _GEN_1174; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1178 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_src2Type : dataBuffer_0_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1179 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_src2Type : _GEN_1178; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1182 = 2'h1 == ringBufferTail ? dataBuffer_1_ctrl_src1Type : dataBuffer_0_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1183 = 2'h2 == ringBufferTail ? dataBuffer_2_ctrl_src1Type : _GEN_1182; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1198 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_crossBoundaryFault : dataBuffer_0_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1199 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_crossBoundaryFault : _GEN_1198; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_1206 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_brIdx : dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [3:0] _GEN_1207 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_brIdx : _GEN_1206; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1214 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_1 : dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1215 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_1 : _GEN_1214; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1222 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_3 : dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1223 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_3 : _GEN_1222; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1230 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_5 : dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1231 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_5 : _GEN_1230; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1238 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_7 : dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1239 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_7 : _GEN_1238; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1246 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_9 : dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1247 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_9 : _GEN_1246; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1254 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_intrVec_11 : dataBuffer_0_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1255 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_intrVec_11 : _GEN_1254; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1262 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_exceptionVec_1 : dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1263 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_exceptionVec_1 : _GEN_1262; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1266 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_exceptionVec_2 : dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1267 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_exceptionVec_2 : _GEN_1266; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1306 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_exceptionVec_12 : dataBuffer_0_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _GEN_1307 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_exceptionVec_12 : _GEN_1306; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_1334 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_pnpc : dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_1335 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_pnpc : _GEN_1334; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_1338 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_pc : dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [38:0] _GEN_1339 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_pc : _GEN_1338; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_1342 = 2'h1 == ringBufferTail ? dataBuffer_1_cf_instr : dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire [63:0] _GEN_1343 = 2'h2 == ringBufferTail ? dataBuffer_2_cf_instr : _GEN_1342; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  wire  _dequeueSize_T = backend_io_in_0_ready & backend_io_in_0_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [1:0] dequeueSize = {{1'd0}, _dequeueSize_T}; // @[src/main/scala/utils/PipelineVector.scala 64:42]
  wire  dequeueFire = dequeueSize > 2'h0; // @[src/main/scala/utils/PipelineVector.scala 65:35]
  wire [1:0] _ringBufferTail_T_1 = ringBufferTail + dequeueSize; // @[src/main/scala/utils/PipelineVector.scala 67:42]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [63:0] dataBuffer_0_cf_instr_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [63:0] dataBuffer_0_cf_instr_t = dataBuffer_0_cf_instr ^ dataBuffer_0_cf_instr_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9135_clock;
  wire  toggle_9135_reset;
  wire [63:0] toggle_9135_valid;
  reg [63:0] toggle_9135_valid_reg;
  reg [38:0] dataBuffer_0_cf_pc_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [38:0] dataBuffer_0_cf_pc_t = dataBuffer_0_cf_pc ^ dataBuffer_0_cf_pc_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9199_clock;
  wire  toggle_9199_reset;
  wire [38:0] toggle_9199_valid;
  reg [38:0] toggle_9199_valid_reg;
  reg [38:0] dataBuffer_0_cf_pnpc_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [38:0] dataBuffer_0_cf_pnpc_t = dataBuffer_0_cf_pnpc ^ dataBuffer_0_cf_pnpc_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9238_clock;
  wire  toggle_9238_reset;
  wire [38:0] toggle_9238_valid;
  reg [38:0] toggle_9238_valid_reg;
  reg  dataBuffer_0_cf_exceptionVec_1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_0_cf_exceptionVec_1_t = dataBuffer_0_cf_exceptionVec_1 ^ dataBuffer_0_cf_exceptionVec_1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9277_clock;
  wire  toggle_9277_reset;
  wire  toggle_9277_valid;
  reg  toggle_9277_valid_reg;
  reg  dataBuffer_0_cf_exceptionVec_2_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_0_cf_exceptionVec_2_t = dataBuffer_0_cf_exceptionVec_2 ^ dataBuffer_0_cf_exceptionVec_2_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9278_clock;
  wire  toggle_9278_reset;
  wire  toggle_9278_valid;
  reg  toggle_9278_valid_reg;
  reg  dataBuffer_0_cf_exceptionVec_12_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_0_cf_exceptionVec_12_t = dataBuffer_0_cf_exceptionVec_12 ^ dataBuffer_0_cf_exceptionVec_12_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9279_clock;
  wire  toggle_9279_reset;
  wire  toggle_9279_valid;
  reg  toggle_9279_valid_reg;
  reg  dataBuffer_0_cf_intrVec_1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_0_cf_intrVec_1_t = dataBuffer_0_cf_intrVec_1 ^ dataBuffer_0_cf_intrVec_1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9280_clock;
  wire  toggle_9280_reset;
  wire  toggle_9280_valid;
  reg  toggle_9280_valid_reg;
  reg  dataBuffer_0_cf_intrVec_3_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_0_cf_intrVec_3_t = dataBuffer_0_cf_intrVec_3 ^ dataBuffer_0_cf_intrVec_3_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9281_clock;
  wire  toggle_9281_reset;
  wire  toggle_9281_valid;
  reg  toggle_9281_valid_reg;
  reg  dataBuffer_0_cf_intrVec_5_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_0_cf_intrVec_5_t = dataBuffer_0_cf_intrVec_5 ^ dataBuffer_0_cf_intrVec_5_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9282_clock;
  wire  toggle_9282_reset;
  wire  toggle_9282_valid;
  reg  toggle_9282_valid_reg;
  reg  dataBuffer_0_cf_intrVec_7_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_0_cf_intrVec_7_t = dataBuffer_0_cf_intrVec_7 ^ dataBuffer_0_cf_intrVec_7_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9283_clock;
  wire  toggle_9283_reset;
  wire  toggle_9283_valid;
  reg  toggle_9283_valid_reg;
  reg  dataBuffer_0_cf_intrVec_9_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_0_cf_intrVec_9_t = dataBuffer_0_cf_intrVec_9 ^ dataBuffer_0_cf_intrVec_9_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9284_clock;
  wire  toggle_9284_reset;
  wire  toggle_9284_valid;
  reg  toggle_9284_valid_reg;
  reg  dataBuffer_0_cf_intrVec_11_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_0_cf_intrVec_11_t = dataBuffer_0_cf_intrVec_11 ^ dataBuffer_0_cf_intrVec_11_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9285_clock;
  wire  toggle_9285_reset;
  wire  toggle_9285_valid;
  reg  toggle_9285_valid_reg;
  reg [3:0] dataBuffer_0_cf_brIdx_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [3:0] dataBuffer_0_cf_brIdx_t = dataBuffer_0_cf_brIdx ^ dataBuffer_0_cf_brIdx_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9286_clock;
  wire  toggle_9286_reset;
  wire [3:0] toggle_9286_valid;
  reg [3:0] toggle_9286_valid_reg;
  reg  dataBuffer_0_cf_crossBoundaryFault_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_0_cf_crossBoundaryFault_t = dataBuffer_0_cf_crossBoundaryFault ^ dataBuffer_0_cf_crossBoundaryFault_p
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9290_clock;
  wire  toggle_9290_reset;
  wire  toggle_9290_valid;
  reg  toggle_9290_valid_reg;
  reg  dataBuffer_0_ctrl_src1Type_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_0_ctrl_src1Type_t = dataBuffer_0_ctrl_src1Type ^ dataBuffer_0_ctrl_src1Type_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9291_clock;
  wire  toggle_9291_reset;
  wire  toggle_9291_valid;
  reg  toggle_9291_valid_reg;
  reg  dataBuffer_0_ctrl_src2Type_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_0_ctrl_src2Type_t = dataBuffer_0_ctrl_src2Type ^ dataBuffer_0_ctrl_src2Type_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9292_clock;
  wire  toggle_9292_reset;
  wire  toggle_9292_valid;
  reg  toggle_9292_valid_reg;
  reg [2:0] dataBuffer_0_ctrl_fuType_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [2:0] dataBuffer_0_ctrl_fuType_t = dataBuffer_0_ctrl_fuType ^ dataBuffer_0_ctrl_fuType_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9293_clock;
  wire  toggle_9293_reset;
  wire [2:0] toggle_9293_valid;
  reg [2:0] toggle_9293_valid_reg;
  reg [6:0] dataBuffer_0_ctrl_fuOpType_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [6:0] dataBuffer_0_ctrl_fuOpType_t = dataBuffer_0_ctrl_fuOpType ^ dataBuffer_0_ctrl_fuOpType_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9296_clock;
  wire  toggle_9296_reset;
  wire [6:0] toggle_9296_valid;
  reg [6:0] toggle_9296_valid_reg;
  reg [4:0] dataBuffer_0_ctrl_rfSrc1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [4:0] dataBuffer_0_ctrl_rfSrc1_t = dataBuffer_0_ctrl_rfSrc1 ^ dataBuffer_0_ctrl_rfSrc1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9303_clock;
  wire  toggle_9303_reset;
  wire [4:0] toggle_9303_valid;
  reg [4:0] toggle_9303_valid_reg;
  reg [4:0] dataBuffer_0_ctrl_rfSrc2_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [4:0] dataBuffer_0_ctrl_rfSrc2_t = dataBuffer_0_ctrl_rfSrc2 ^ dataBuffer_0_ctrl_rfSrc2_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9308_clock;
  wire  toggle_9308_reset;
  wire [4:0] toggle_9308_valid;
  reg [4:0] toggle_9308_valid_reg;
  reg  dataBuffer_0_ctrl_rfWen_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_0_ctrl_rfWen_t = dataBuffer_0_ctrl_rfWen ^ dataBuffer_0_ctrl_rfWen_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9313_clock;
  wire  toggle_9313_reset;
  wire  toggle_9313_valid;
  reg  toggle_9313_valid_reg;
  reg [4:0] dataBuffer_0_ctrl_rfDest_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [4:0] dataBuffer_0_ctrl_rfDest_t = dataBuffer_0_ctrl_rfDest ^ dataBuffer_0_ctrl_rfDest_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9314_clock;
  wire  toggle_9314_reset;
  wire [4:0] toggle_9314_valid;
  reg [4:0] toggle_9314_valid_reg;
  reg  dataBuffer_0_ctrl_isNutCoreTrap_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_0_ctrl_isNutCoreTrap_t = dataBuffer_0_ctrl_isNutCoreTrap ^ dataBuffer_0_ctrl_isNutCoreTrap_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9319_clock;
  wire  toggle_9319_reset;
  wire  toggle_9319_valid;
  reg  toggle_9319_valid_reg;
  reg [63:0] dataBuffer_0_data_imm_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [63:0] dataBuffer_0_data_imm_t = dataBuffer_0_data_imm ^ dataBuffer_0_data_imm_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9320_clock;
  wire  toggle_9320_reset;
  wire [63:0] toggle_9320_valid;
  reg [63:0] toggle_9320_valid_reg;
  reg [63:0] dataBuffer_1_cf_instr_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [63:0] dataBuffer_1_cf_instr_t = dataBuffer_1_cf_instr ^ dataBuffer_1_cf_instr_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9384_clock;
  wire  toggle_9384_reset;
  wire [63:0] toggle_9384_valid;
  reg [63:0] toggle_9384_valid_reg;
  reg [38:0] dataBuffer_1_cf_pc_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [38:0] dataBuffer_1_cf_pc_t = dataBuffer_1_cf_pc ^ dataBuffer_1_cf_pc_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9448_clock;
  wire  toggle_9448_reset;
  wire [38:0] toggle_9448_valid;
  reg [38:0] toggle_9448_valid_reg;
  reg [38:0] dataBuffer_1_cf_pnpc_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [38:0] dataBuffer_1_cf_pnpc_t = dataBuffer_1_cf_pnpc ^ dataBuffer_1_cf_pnpc_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9487_clock;
  wire  toggle_9487_reset;
  wire [38:0] toggle_9487_valid;
  reg [38:0] toggle_9487_valid_reg;
  reg  dataBuffer_1_cf_exceptionVec_1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_1_cf_exceptionVec_1_t = dataBuffer_1_cf_exceptionVec_1 ^ dataBuffer_1_cf_exceptionVec_1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9526_clock;
  wire  toggle_9526_reset;
  wire  toggle_9526_valid;
  reg  toggle_9526_valid_reg;
  reg  dataBuffer_1_cf_exceptionVec_2_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_1_cf_exceptionVec_2_t = dataBuffer_1_cf_exceptionVec_2 ^ dataBuffer_1_cf_exceptionVec_2_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9527_clock;
  wire  toggle_9527_reset;
  wire  toggle_9527_valid;
  reg  toggle_9527_valid_reg;
  reg  dataBuffer_1_cf_exceptionVec_12_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_1_cf_exceptionVec_12_t = dataBuffer_1_cf_exceptionVec_12 ^ dataBuffer_1_cf_exceptionVec_12_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9528_clock;
  wire  toggle_9528_reset;
  wire  toggle_9528_valid;
  reg  toggle_9528_valid_reg;
  reg  dataBuffer_1_cf_intrVec_1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_1_cf_intrVec_1_t = dataBuffer_1_cf_intrVec_1 ^ dataBuffer_1_cf_intrVec_1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9529_clock;
  wire  toggle_9529_reset;
  wire  toggle_9529_valid;
  reg  toggle_9529_valid_reg;
  reg  dataBuffer_1_cf_intrVec_3_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_1_cf_intrVec_3_t = dataBuffer_1_cf_intrVec_3 ^ dataBuffer_1_cf_intrVec_3_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9530_clock;
  wire  toggle_9530_reset;
  wire  toggle_9530_valid;
  reg  toggle_9530_valid_reg;
  reg  dataBuffer_1_cf_intrVec_5_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_1_cf_intrVec_5_t = dataBuffer_1_cf_intrVec_5 ^ dataBuffer_1_cf_intrVec_5_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9531_clock;
  wire  toggle_9531_reset;
  wire  toggle_9531_valid;
  reg  toggle_9531_valid_reg;
  reg  dataBuffer_1_cf_intrVec_7_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_1_cf_intrVec_7_t = dataBuffer_1_cf_intrVec_7 ^ dataBuffer_1_cf_intrVec_7_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9532_clock;
  wire  toggle_9532_reset;
  wire  toggle_9532_valid;
  reg  toggle_9532_valid_reg;
  reg  dataBuffer_1_cf_intrVec_9_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_1_cf_intrVec_9_t = dataBuffer_1_cf_intrVec_9 ^ dataBuffer_1_cf_intrVec_9_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9533_clock;
  wire  toggle_9533_reset;
  wire  toggle_9533_valid;
  reg  toggle_9533_valid_reg;
  reg  dataBuffer_1_cf_intrVec_11_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_1_cf_intrVec_11_t = dataBuffer_1_cf_intrVec_11 ^ dataBuffer_1_cf_intrVec_11_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9534_clock;
  wire  toggle_9534_reset;
  wire  toggle_9534_valid;
  reg  toggle_9534_valid_reg;
  reg [3:0] dataBuffer_1_cf_brIdx_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [3:0] dataBuffer_1_cf_brIdx_t = dataBuffer_1_cf_brIdx ^ dataBuffer_1_cf_brIdx_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9535_clock;
  wire  toggle_9535_reset;
  wire [3:0] toggle_9535_valid;
  reg [3:0] toggle_9535_valid_reg;
  reg  dataBuffer_1_cf_crossBoundaryFault_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_1_cf_crossBoundaryFault_t = dataBuffer_1_cf_crossBoundaryFault ^ dataBuffer_1_cf_crossBoundaryFault_p
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9539_clock;
  wire  toggle_9539_reset;
  wire  toggle_9539_valid;
  reg  toggle_9539_valid_reg;
  reg  dataBuffer_1_ctrl_src1Type_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_1_ctrl_src1Type_t = dataBuffer_1_ctrl_src1Type ^ dataBuffer_1_ctrl_src1Type_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9540_clock;
  wire  toggle_9540_reset;
  wire  toggle_9540_valid;
  reg  toggle_9540_valid_reg;
  reg  dataBuffer_1_ctrl_src2Type_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_1_ctrl_src2Type_t = dataBuffer_1_ctrl_src2Type ^ dataBuffer_1_ctrl_src2Type_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9541_clock;
  wire  toggle_9541_reset;
  wire  toggle_9541_valid;
  reg  toggle_9541_valid_reg;
  reg [2:0] dataBuffer_1_ctrl_fuType_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [2:0] dataBuffer_1_ctrl_fuType_t = dataBuffer_1_ctrl_fuType ^ dataBuffer_1_ctrl_fuType_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9542_clock;
  wire  toggle_9542_reset;
  wire [2:0] toggle_9542_valid;
  reg [2:0] toggle_9542_valid_reg;
  reg [6:0] dataBuffer_1_ctrl_fuOpType_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [6:0] dataBuffer_1_ctrl_fuOpType_t = dataBuffer_1_ctrl_fuOpType ^ dataBuffer_1_ctrl_fuOpType_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9545_clock;
  wire  toggle_9545_reset;
  wire [6:0] toggle_9545_valid;
  reg [6:0] toggle_9545_valid_reg;
  reg [4:0] dataBuffer_1_ctrl_rfSrc1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [4:0] dataBuffer_1_ctrl_rfSrc1_t = dataBuffer_1_ctrl_rfSrc1 ^ dataBuffer_1_ctrl_rfSrc1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9552_clock;
  wire  toggle_9552_reset;
  wire [4:0] toggle_9552_valid;
  reg [4:0] toggle_9552_valid_reg;
  reg [4:0] dataBuffer_1_ctrl_rfSrc2_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [4:0] dataBuffer_1_ctrl_rfSrc2_t = dataBuffer_1_ctrl_rfSrc2 ^ dataBuffer_1_ctrl_rfSrc2_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9557_clock;
  wire  toggle_9557_reset;
  wire [4:0] toggle_9557_valid;
  reg [4:0] toggle_9557_valid_reg;
  reg  dataBuffer_1_ctrl_rfWen_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_1_ctrl_rfWen_t = dataBuffer_1_ctrl_rfWen ^ dataBuffer_1_ctrl_rfWen_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9562_clock;
  wire  toggle_9562_reset;
  wire  toggle_9562_valid;
  reg  toggle_9562_valid_reg;
  reg [4:0] dataBuffer_1_ctrl_rfDest_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [4:0] dataBuffer_1_ctrl_rfDest_t = dataBuffer_1_ctrl_rfDest ^ dataBuffer_1_ctrl_rfDest_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9563_clock;
  wire  toggle_9563_reset;
  wire [4:0] toggle_9563_valid;
  reg [4:0] toggle_9563_valid_reg;
  reg  dataBuffer_1_ctrl_isNutCoreTrap_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_1_ctrl_isNutCoreTrap_t = dataBuffer_1_ctrl_isNutCoreTrap ^ dataBuffer_1_ctrl_isNutCoreTrap_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9568_clock;
  wire  toggle_9568_reset;
  wire  toggle_9568_valid;
  reg  toggle_9568_valid_reg;
  reg [63:0] dataBuffer_1_data_imm_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [63:0] dataBuffer_1_data_imm_t = dataBuffer_1_data_imm ^ dataBuffer_1_data_imm_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9569_clock;
  wire  toggle_9569_reset;
  wire [63:0] toggle_9569_valid;
  reg [63:0] toggle_9569_valid_reg;
  reg [63:0] dataBuffer_2_cf_instr_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [63:0] dataBuffer_2_cf_instr_t = dataBuffer_2_cf_instr ^ dataBuffer_2_cf_instr_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9633_clock;
  wire  toggle_9633_reset;
  wire [63:0] toggle_9633_valid;
  reg [63:0] toggle_9633_valid_reg;
  reg [38:0] dataBuffer_2_cf_pc_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [38:0] dataBuffer_2_cf_pc_t = dataBuffer_2_cf_pc ^ dataBuffer_2_cf_pc_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9697_clock;
  wire  toggle_9697_reset;
  wire [38:0] toggle_9697_valid;
  reg [38:0] toggle_9697_valid_reg;
  reg [38:0] dataBuffer_2_cf_pnpc_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [38:0] dataBuffer_2_cf_pnpc_t = dataBuffer_2_cf_pnpc ^ dataBuffer_2_cf_pnpc_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9736_clock;
  wire  toggle_9736_reset;
  wire [38:0] toggle_9736_valid;
  reg [38:0] toggle_9736_valid_reg;
  reg  dataBuffer_2_cf_exceptionVec_1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_2_cf_exceptionVec_1_t = dataBuffer_2_cf_exceptionVec_1 ^ dataBuffer_2_cf_exceptionVec_1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9775_clock;
  wire  toggle_9775_reset;
  wire  toggle_9775_valid;
  reg  toggle_9775_valid_reg;
  reg  dataBuffer_2_cf_exceptionVec_2_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_2_cf_exceptionVec_2_t = dataBuffer_2_cf_exceptionVec_2 ^ dataBuffer_2_cf_exceptionVec_2_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9776_clock;
  wire  toggle_9776_reset;
  wire  toggle_9776_valid;
  reg  toggle_9776_valid_reg;
  reg  dataBuffer_2_cf_exceptionVec_12_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_2_cf_exceptionVec_12_t = dataBuffer_2_cf_exceptionVec_12 ^ dataBuffer_2_cf_exceptionVec_12_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9777_clock;
  wire  toggle_9777_reset;
  wire  toggle_9777_valid;
  reg  toggle_9777_valid_reg;
  reg  dataBuffer_2_cf_intrVec_1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_2_cf_intrVec_1_t = dataBuffer_2_cf_intrVec_1 ^ dataBuffer_2_cf_intrVec_1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9778_clock;
  wire  toggle_9778_reset;
  wire  toggle_9778_valid;
  reg  toggle_9778_valid_reg;
  reg  dataBuffer_2_cf_intrVec_3_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_2_cf_intrVec_3_t = dataBuffer_2_cf_intrVec_3 ^ dataBuffer_2_cf_intrVec_3_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9779_clock;
  wire  toggle_9779_reset;
  wire  toggle_9779_valid;
  reg  toggle_9779_valid_reg;
  reg  dataBuffer_2_cf_intrVec_5_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_2_cf_intrVec_5_t = dataBuffer_2_cf_intrVec_5 ^ dataBuffer_2_cf_intrVec_5_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9780_clock;
  wire  toggle_9780_reset;
  wire  toggle_9780_valid;
  reg  toggle_9780_valid_reg;
  reg  dataBuffer_2_cf_intrVec_7_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_2_cf_intrVec_7_t = dataBuffer_2_cf_intrVec_7 ^ dataBuffer_2_cf_intrVec_7_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9781_clock;
  wire  toggle_9781_reset;
  wire  toggle_9781_valid;
  reg  toggle_9781_valid_reg;
  reg  dataBuffer_2_cf_intrVec_9_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_2_cf_intrVec_9_t = dataBuffer_2_cf_intrVec_9 ^ dataBuffer_2_cf_intrVec_9_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9782_clock;
  wire  toggle_9782_reset;
  wire  toggle_9782_valid;
  reg  toggle_9782_valid_reg;
  reg  dataBuffer_2_cf_intrVec_11_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_2_cf_intrVec_11_t = dataBuffer_2_cf_intrVec_11 ^ dataBuffer_2_cf_intrVec_11_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9783_clock;
  wire  toggle_9783_reset;
  wire  toggle_9783_valid;
  reg  toggle_9783_valid_reg;
  reg [3:0] dataBuffer_2_cf_brIdx_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [3:0] dataBuffer_2_cf_brIdx_t = dataBuffer_2_cf_brIdx ^ dataBuffer_2_cf_brIdx_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9784_clock;
  wire  toggle_9784_reset;
  wire [3:0] toggle_9784_valid;
  reg [3:0] toggle_9784_valid_reg;
  reg  dataBuffer_2_cf_crossBoundaryFault_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_2_cf_crossBoundaryFault_t = dataBuffer_2_cf_crossBoundaryFault ^ dataBuffer_2_cf_crossBoundaryFault_p
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9788_clock;
  wire  toggle_9788_reset;
  wire  toggle_9788_valid;
  reg  toggle_9788_valid_reg;
  reg  dataBuffer_2_ctrl_src1Type_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_2_ctrl_src1Type_t = dataBuffer_2_ctrl_src1Type ^ dataBuffer_2_ctrl_src1Type_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9789_clock;
  wire  toggle_9789_reset;
  wire  toggle_9789_valid;
  reg  toggle_9789_valid_reg;
  reg  dataBuffer_2_ctrl_src2Type_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_2_ctrl_src2Type_t = dataBuffer_2_ctrl_src2Type ^ dataBuffer_2_ctrl_src2Type_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9790_clock;
  wire  toggle_9790_reset;
  wire  toggle_9790_valid;
  reg  toggle_9790_valid_reg;
  reg [2:0] dataBuffer_2_ctrl_fuType_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [2:0] dataBuffer_2_ctrl_fuType_t = dataBuffer_2_ctrl_fuType ^ dataBuffer_2_ctrl_fuType_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9791_clock;
  wire  toggle_9791_reset;
  wire [2:0] toggle_9791_valid;
  reg [2:0] toggle_9791_valid_reg;
  reg [6:0] dataBuffer_2_ctrl_fuOpType_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [6:0] dataBuffer_2_ctrl_fuOpType_t = dataBuffer_2_ctrl_fuOpType ^ dataBuffer_2_ctrl_fuOpType_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9794_clock;
  wire  toggle_9794_reset;
  wire [6:0] toggle_9794_valid;
  reg [6:0] toggle_9794_valid_reg;
  reg [4:0] dataBuffer_2_ctrl_rfSrc1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [4:0] dataBuffer_2_ctrl_rfSrc1_t = dataBuffer_2_ctrl_rfSrc1 ^ dataBuffer_2_ctrl_rfSrc1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9801_clock;
  wire  toggle_9801_reset;
  wire [4:0] toggle_9801_valid;
  reg [4:0] toggle_9801_valid_reg;
  reg [4:0] dataBuffer_2_ctrl_rfSrc2_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [4:0] dataBuffer_2_ctrl_rfSrc2_t = dataBuffer_2_ctrl_rfSrc2 ^ dataBuffer_2_ctrl_rfSrc2_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9806_clock;
  wire  toggle_9806_reset;
  wire [4:0] toggle_9806_valid;
  reg [4:0] toggle_9806_valid_reg;
  reg  dataBuffer_2_ctrl_rfWen_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_2_ctrl_rfWen_t = dataBuffer_2_ctrl_rfWen ^ dataBuffer_2_ctrl_rfWen_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9811_clock;
  wire  toggle_9811_reset;
  wire  toggle_9811_valid;
  reg  toggle_9811_valid_reg;
  reg [4:0] dataBuffer_2_ctrl_rfDest_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [4:0] dataBuffer_2_ctrl_rfDest_t = dataBuffer_2_ctrl_rfDest ^ dataBuffer_2_ctrl_rfDest_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9812_clock;
  wire  toggle_9812_reset;
  wire [4:0] toggle_9812_valid;
  reg [4:0] toggle_9812_valid_reg;
  reg  dataBuffer_2_ctrl_isNutCoreTrap_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_2_ctrl_isNutCoreTrap_t = dataBuffer_2_ctrl_isNutCoreTrap ^ dataBuffer_2_ctrl_isNutCoreTrap_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9817_clock;
  wire  toggle_9817_reset;
  wire  toggle_9817_valid;
  reg  toggle_9817_valid_reg;
  reg [63:0] dataBuffer_2_data_imm_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [63:0] dataBuffer_2_data_imm_t = dataBuffer_2_data_imm ^ dataBuffer_2_data_imm_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9818_clock;
  wire  toggle_9818_reset;
  wire [63:0] toggle_9818_valid;
  reg [63:0] toggle_9818_valid_reg;
  reg [63:0] dataBuffer_3_cf_instr_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [63:0] dataBuffer_3_cf_instr_t = dataBuffer_3_cf_instr ^ dataBuffer_3_cf_instr_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9882_clock;
  wire  toggle_9882_reset;
  wire [63:0] toggle_9882_valid;
  reg [63:0] toggle_9882_valid_reg;
  reg [38:0] dataBuffer_3_cf_pc_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [38:0] dataBuffer_3_cf_pc_t = dataBuffer_3_cf_pc ^ dataBuffer_3_cf_pc_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9946_clock;
  wire  toggle_9946_reset;
  wire [38:0] toggle_9946_valid;
  reg [38:0] toggle_9946_valid_reg;
  reg [38:0] dataBuffer_3_cf_pnpc_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [38:0] dataBuffer_3_cf_pnpc_t = dataBuffer_3_cf_pnpc ^ dataBuffer_3_cf_pnpc_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_9985_clock;
  wire  toggle_9985_reset;
  wire [38:0] toggle_9985_valid;
  reg [38:0] toggle_9985_valid_reg;
  reg  dataBuffer_3_cf_exceptionVec_1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_3_cf_exceptionVec_1_t = dataBuffer_3_cf_exceptionVec_1 ^ dataBuffer_3_cf_exceptionVec_1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10024_clock;
  wire  toggle_10024_reset;
  wire  toggle_10024_valid;
  reg  toggle_10024_valid_reg;
  reg  dataBuffer_3_cf_exceptionVec_2_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_3_cf_exceptionVec_2_t = dataBuffer_3_cf_exceptionVec_2 ^ dataBuffer_3_cf_exceptionVec_2_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10025_clock;
  wire  toggle_10025_reset;
  wire  toggle_10025_valid;
  reg  toggle_10025_valid_reg;
  reg  dataBuffer_3_cf_exceptionVec_12_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_3_cf_exceptionVec_12_t = dataBuffer_3_cf_exceptionVec_12 ^ dataBuffer_3_cf_exceptionVec_12_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10026_clock;
  wire  toggle_10026_reset;
  wire  toggle_10026_valid;
  reg  toggle_10026_valid_reg;
  reg  dataBuffer_3_cf_intrVec_1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_3_cf_intrVec_1_t = dataBuffer_3_cf_intrVec_1 ^ dataBuffer_3_cf_intrVec_1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10027_clock;
  wire  toggle_10027_reset;
  wire  toggle_10027_valid;
  reg  toggle_10027_valid_reg;
  reg  dataBuffer_3_cf_intrVec_3_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_3_cf_intrVec_3_t = dataBuffer_3_cf_intrVec_3 ^ dataBuffer_3_cf_intrVec_3_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10028_clock;
  wire  toggle_10028_reset;
  wire  toggle_10028_valid;
  reg  toggle_10028_valid_reg;
  reg  dataBuffer_3_cf_intrVec_5_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_3_cf_intrVec_5_t = dataBuffer_3_cf_intrVec_5 ^ dataBuffer_3_cf_intrVec_5_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10029_clock;
  wire  toggle_10029_reset;
  wire  toggle_10029_valid;
  reg  toggle_10029_valid_reg;
  reg  dataBuffer_3_cf_intrVec_7_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_3_cf_intrVec_7_t = dataBuffer_3_cf_intrVec_7 ^ dataBuffer_3_cf_intrVec_7_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10030_clock;
  wire  toggle_10030_reset;
  wire  toggle_10030_valid;
  reg  toggle_10030_valid_reg;
  reg  dataBuffer_3_cf_intrVec_9_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_3_cf_intrVec_9_t = dataBuffer_3_cf_intrVec_9 ^ dataBuffer_3_cf_intrVec_9_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10031_clock;
  wire  toggle_10031_reset;
  wire  toggle_10031_valid;
  reg  toggle_10031_valid_reg;
  reg  dataBuffer_3_cf_intrVec_11_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_3_cf_intrVec_11_t = dataBuffer_3_cf_intrVec_11 ^ dataBuffer_3_cf_intrVec_11_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10032_clock;
  wire  toggle_10032_reset;
  wire  toggle_10032_valid;
  reg  toggle_10032_valid_reg;
  reg [3:0] dataBuffer_3_cf_brIdx_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [3:0] dataBuffer_3_cf_brIdx_t = dataBuffer_3_cf_brIdx ^ dataBuffer_3_cf_brIdx_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10033_clock;
  wire  toggle_10033_reset;
  wire [3:0] toggle_10033_valid;
  reg [3:0] toggle_10033_valid_reg;
  reg  dataBuffer_3_cf_crossBoundaryFault_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_3_cf_crossBoundaryFault_t = dataBuffer_3_cf_crossBoundaryFault ^ dataBuffer_3_cf_crossBoundaryFault_p
    ; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10037_clock;
  wire  toggle_10037_reset;
  wire  toggle_10037_valid;
  reg  toggle_10037_valid_reg;
  reg  dataBuffer_3_ctrl_src1Type_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_3_ctrl_src1Type_t = dataBuffer_3_ctrl_src1Type ^ dataBuffer_3_ctrl_src1Type_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10038_clock;
  wire  toggle_10038_reset;
  wire  toggle_10038_valid;
  reg  toggle_10038_valid_reg;
  reg  dataBuffer_3_ctrl_src2Type_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_3_ctrl_src2Type_t = dataBuffer_3_ctrl_src2Type ^ dataBuffer_3_ctrl_src2Type_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10039_clock;
  wire  toggle_10039_reset;
  wire  toggle_10039_valid;
  reg  toggle_10039_valid_reg;
  reg [2:0] dataBuffer_3_ctrl_fuType_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [2:0] dataBuffer_3_ctrl_fuType_t = dataBuffer_3_ctrl_fuType ^ dataBuffer_3_ctrl_fuType_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10040_clock;
  wire  toggle_10040_reset;
  wire [2:0] toggle_10040_valid;
  reg [2:0] toggle_10040_valid_reg;
  reg [6:0] dataBuffer_3_ctrl_fuOpType_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [6:0] dataBuffer_3_ctrl_fuOpType_t = dataBuffer_3_ctrl_fuOpType ^ dataBuffer_3_ctrl_fuOpType_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10043_clock;
  wire  toggle_10043_reset;
  wire [6:0] toggle_10043_valid;
  reg [6:0] toggle_10043_valid_reg;
  reg [4:0] dataBuffer_3_ctrl_rfSrc1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [4:0] dataBuffer_3_ctrl_rfSrc1_t = dataBuffer_3_ctrl_rfSrc1 ^ dataBuffer_3_ctrl_rfSrc1_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10050_clock;
  wire  toggle_10050_reset;
  wire [4:0] toggle_10050_valid;
  reg [4:0] toggle_10050_valid_reg;
  reg [4:0] dataBuffer_3_ctrl_rfSrc2_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [4:0] dataBuffer_3_ctrl_rfSrc2_t = dataBuffer_3_ctrl_rfSrc2 ^ dataBuffer_3_ctrl_rfSrc2_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10055_clock;
  wire  toggle_10055_reset;
  wire [4:0] toggle_10055_valid;
  reg [4:0] toggle_10055_valid_reg;
  reg  dataBuffer_3_ctrl_rfWen_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_3_ctrl_rfWen_t = dataBuffer_3_ctrl_rfWen ^ dataBuffer_3_ctrl_rfWen_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10060_clock;
  wire  toggle_10060_reset;
  wire  toggle_10060_valid;
  reg  toggle_10060_valid_reg;
  reg [4:0] dataBuffer_3_ctrl_rfDest_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [4:0] dataBuffer_3_ctrl_rfDest_t = dataBuffer_3_ctrl_rfDest ^ dataBuffer_3_ctrl_rfDest_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10061_clock;
  wire  toggle_10061_reset;
  wire [4:0] toggle_10061_valid;
  reg [4:0] toggle_10061_valid_reg;
  reg  dataBuffer_3_ctrl_isNutCoreTrap_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  dataBuffer_3_ctrl_isNutCoreTrap_t = dataBuffer_3_ctrl_isNutCoreTrap ^ dataBuffer_3_ctrl_isNutCoreTrap_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10066_clock;
  wire  toggle_10066_reset;
  wire  toggle_10066_valid;
  reg  toggle_10066_valid_reg;
  reg [63:0] dataBuffer_3_data_imm_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire [63:0] dataBuffer_3_data_imm_t = dataBuffer_3_data_imm ^ dataBuffer_3_data_imm_p; // @[src/main/scala/utils/PipelineVector.scala 29:29]
  wire  toggle_10067_clock;
  wire  toggle_10067_reset;
  wire [63:0] toggle_10067_valid;
  reg [63:0] toggle_10067_valid_reg;
  reg [1:0] ringBufferHead_p; // @[src/main/scala/utils/PipelineVector.scala 30:33]
  wire [1:0] ringBufferHead_t = ringBufferHead ^ ringBufferHead_p; // @[src/main/scala/utils/PipelineVector.scala 30:33]
  wire  toggle_10131_clock;
  wire  toggle_10131_reset;
  wire [1:0] toggle_10131_valid;
  reg [1:0] toggle_10131_valid_reg;
  reg [1:0] ringBufferTail_p; // @[src/main/scala/utils/PipelineVector.scala 31:33]
  wire [1:0] ringBufferTail_t = ringBufferTail ^ ringBufferTail_p; // @[src/main/scala/utils/PipelineVector.scala 31:33]
  wire  toggle_10133_clock;
  wire  toggle_10133_reset;
  wire [1:0] toggle_10133_valid;
  reg [1:0] toggle_10133_valid_reg;
  Frontend_inorder frontend ( // @[src/main/scala/nutcore/NutCore.scala 131:34]
    .clock(frontend_clock),
    .reset(frontend_reset),
    .io_imem_req_ready(frontend_io_imem_req_ready),
    .io_imem_req_valid(frontend_io_imem_req_valid),
    .io_imem_req_bits_addr(frontend_io_imem_req_bits_addr),
    .io_imem_req_bits_user(frontend_io_imem_req_bits_user),
    .io_imem_resp_ready(frontend_io_imem_resp_ready),
    .io_imem_resp_valid(frontend_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(frontend_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(frontend_io_imem_resp_bits_user),
    .io_out_0_ready(frontend_io_out_0_ready),
    .io_out_0_valid(frontend_io_out_0_valid),
    .io_out_0_bits_cf_instr(frontend_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(frontend_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(frontend_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(frontend_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(frontend_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(frontend_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_intrVec_1(frontend_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_3(frontend_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_5(frontend_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_7(frontend_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_9(frontend_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_11(frontend_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(frontend_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_cf_crossBoundaryFault(frontend_io_out_0_bits_cf_crossBoundaryFault),
    .io_out_0_bits_ctrl_src1Type(frontend_io_out_0_bits_ctrl_src1Type),
    .io_out_0_bits_ctrl_src2Type(frontend_io_out_0_bits_ctrl_src2Type),
    .io_out_0_bits_ctrl_fuType(frontend_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(frontend_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfSrc1(frontend_io_out_0_bits_ctrl_rfSrc1),
    .io_out_0_bits_ctrl_rfSrc2(frontend_io_out_0_bits_ctrl_rfSrc2),
    .io_out_0_bits_ctrl_rfWen(frontend_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(frontend_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_ctrl_isNutCoreTrap(frontend_io_out_0_bits_ctrl_isNutCoreTrap),
    .io_out_0_bits_data_imm(frontend_io_out_0_bits_data_imm),
    .io_flushVec(frontend_io_flushVec),
    .io_redirect_target(frontend_io_redirect_target),
    .io_redirect_valid(frontend_io_redirect_valid),
    .io_iaf(frontend_io_iaf),
    .io_sfence_vma_invalid(frontend_io_sfence_vma_invalid),
    .io_wfi_invalid(frontend_io_wfi_invalid),
    .REG_valid(frontend_REG_valid),
    .REG_pc(frontend_REG_pc),
    .REG_isMissPredict(frontend_REG_isMissPredict),
    .REG_actualTarget(frontend_REG_actualTarget),
    .REG_fuOpType(frontend_REG_fuOpType),
    .REG_btbType(frontend_REG_btbType),
    .REG_isRVC(frontend_REG_isRVC),
    .isWFI(frontend_isWFI),
    .flushICache(frontend_flushICache),
    .flushTLB(frontend_flushTLB),
    .intrVecIDU(frontend_intrVecIDU)
  );
  Backend_inorder backend ( // @[src/main/scala/nutcore/NutCore.scala 174:25]
    .clock(backend_clock),
    .reset(backend_reset),
    .io_in_0_ready(backend_io_in_0_ready),
    .io_in_0_valid(backend_io_in_0_valid),
    .io_in_0_bits_cf_instr(backend_io_in_0_bits_cf_instr),
    .io_in_0_bits_cf_pc(backend_io_in_0_bits_cf_pc),
    .io_in_0_bits_cf_pnpc(backend_io_in_0_bits_cf_pnpc),
    .io_in_0_bits_cf_exceptionVec_1(backend_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(backend_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_exceptionVec_12(backend_io_in_0_bits_cf_exceptionVec_12),
    .io_in_0_bits_cf_intrVec_1(backend_io_in_0_bits_cf_intrVec_1),
    .io_in_0_bits_cf_intrVec_3(backend_io_in_0_bits_cf_intrVec_3),
    .io_in_0_bits_cf_intrVec_5(backend_io_in_0_bits_cf_intrVec_5),
    .io_in_0_bits_cf_intrVec_7(backend_io_in_0_bits_cf_intrVec_7),
    .io_in_0_bits_cf_intrVec_9(backend_io_in_0_bits_cf_intrVec_9),
    .io_in_0_bits_cf_intrVec_11(backend_io_in_0_bits_cf_intrVec_11),
    .io_in_0_bits_cf_brIdx(backend_io_in_0_bits_cf_brIdx),
    .io_in_0_bits_cf_crossBoundaryFault(backend_io_in_0_bits_cf_crossBoundaryFault),
    .io_in_0_bits_ctrl_src1Type(backend_io_in_0_bits_ctrl_src1Type),
    .io_in_0_bits_ctrl_src2Type(backend_io_in_0_bits_ctrl_src2Type),
    .io_in_0_bits_ctrl_fuType(backend_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(backend_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_rfSrc1(backend_io_in_0_bits_ctrl_rfSrc1),
    .io_in_0_bits_ctrl_rfSrc2(backend_io_in_0_bits_ctrl_rfSrc2),
    .io_in_0_bits_ctrl_rfWen(backend_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_rfDest(backend_io_in_0_bits_ctrl_rfDest),
    .io_in_0_bits_ctrl_isNutCoreTrap(backend_io_in_0_bits_ctrl_isNutCoreTrap),
    .io_in_0_bits_data_imm(backend_io_in_0_bits_data_imm),
    .io_flush(backend_io_flush),
    .io_dmem_req_ready(backend_io_dmem_req_ready),
    .io_dmem_req_valid(backend_io_dmem_req_valid),
    .io_dmem_req_bits_addr(backend_io_dmem_req_bits_addr),
    .io_dmem_req_bits_size(backend_io_dmem_req_bits_size),
    .io_dmem_req_bits_cmd(backend_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_wmask(backend_io_dmem_req_bits_wmask),
    .io_dmem_req_bits_wdata(backend_io_dmem_req_bits_wdata),
    .io_dmem_resp_valid(backend_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(backend_io_dmem_resp_bits_rdata),
    .io_memMMU_imem_priviledgeMode(backend_io_memMMU_imem_priviledgeMode),
    .io_memMMU_dmem_priviledgeMode(backend_io_memMMU_dmem_priviledgeMode),
    .io_memMMU_dmem_status_sum(backend_io_memMMU_dmem_status_sum),
    .io_memMMU_dmem_status_mxr(backend_io_memMMU_dmem_status_mxr),
    .io_memMMU_dmem_loadPF(backend_io_memMMU_dmem_loadPF),
    .io_memMMU_dmem_storePF(backend_io_memMMU_dmem_storePF),
    .io_memMMU_dmem_laf(backend_io_memMMU_dmem_laf),
    .io_memMMU_dmem_saf(backend_io_memMMU_dmem_saf),
    .io_sfence_vma_invalid(backend_io_sfence_vma_invalid),
    .io_wfi_invalid(backend_io_wfi_invalid),
    .io_redirect_target(backend_io_redirect_target),
    .io_redirect_valid(backend_io_redirect_valid),
    .lr(backend_lr),
    .io_extra_meip_0(backend_io_extra_meip_0),
    .scInflight(backend_scInflight),
    .REG_valid(backend_REG_valid),
    .REG_pc(backend_REG_pc),
    .REG_isMissPredict(backend_REG_isMissPredict),
    .REG_actualTarget(backend_REG_actualTarget),
    .REG_fuOpType(backend_REG_fuOpType),
    .REG_btbType(backend_REG_btbType),
    .REG_isRVC(backend_REG_isRVC),
    .amoReq(backend_amoReq),
    .lrAddr(backend_lrAddr),
    .paddr(backend_paddr),
    .satp(backend_satp),
    ._T_12(backend__T_12),
    .scIsSuccess(backend_scIsSuccess),
    .io_extra_mtip(backend_io_extra_mtip),
    .flushICache(backend_flushICache),
    .vmEnable(backend_vmEnable),
    .flushTLB(backend_flushTLB),
    .intrVecIDU(backend_intrVecIDU),
    .tlbFinish(backend_tlbFinish),
    .ismmio(backend_ismmio),
    ._T_13_0(backend__T_13_0),
    .io_extra_msip(backend_io_extra_msip)
  );
  SimpleBusCrossbarNto1 mmioXbar ( // @[src/main/scala/nutcore/NutCore.scala 178:26]
    .clock(mmioXbar_clock),
    .reset(mmioXbar_reset),
    .io_in_0_req_ready(mmioXbar_io_in_0_req_ready),
    .io_in_0_req_valid(mmioXbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(mmioXbar_io_in_0_req_bits_addr),
    .io_in_0_resp_valid(mmioXbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_rdata(mmioXbar_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(mmioXbar_io_in_1_req_ready),
    .io_in_1_req_valid(mmioXbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(mmioXbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_cmd(mmioXbar_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(mmioXbar_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(mmioXbar_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(mmioXbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(mmioXbar_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(mmioXbar_io_in_1_resp_bits_rdata),
    .io_out_req_ready(mmioXbar_io_out_req_ready),
    .io_out_req_valid(mmioXbar_io_out_req_valid),
    .io_out_req_bits_addr(mmioXbar_io_out_req_bits_addr),
    .io_out_req_bits_cmd(mmioXbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(mmioXbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(mmioXbar_io_out_req_bits_wdata),
    .io_out_resp_ready(mmioXbar_io_out_resp_ready),
    .io_out_resp_valid(mmioXbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(mmioXbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(mmioXbar_io_out_resp_bits_rdata)
  );
  SimpleBusCrossbarNto1_1 dmemXbar ( // @[src/main/scala/nutcore/NutCore.scala 179:26]
    .clock(dmemXbar_clock),
    .reset(dmemXbar_reset),
    .io_in_0_req_ready(dmemXbar_io_in_0_req_ready),
    .io_in_0_req_valid(dmemXbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(dmemXbar_io_in_0_req_bits_addr),
    .io_in_0_req_bits_size(dmemXbar_io_in_0_req_bits_size),
    .io_in_0_req_bits_cmd(dmemXbar_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(dmemXbar_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(dmemXbar_io_in_0_req_bits_wdata),
    .io_in_0_resp_valid(dmemXbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_rdata(dmemXbar_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(dmemXbar_io_in_1_req_ready),
    .io_in_1_req_valid(dmemXbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(dmemXbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_cmd(dmemXbar_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wdata(dmemXbar_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(dmemXbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_rdata(dmemXbar_io_in_1_resp_bits_rdata),
    .io_in_2_req_ready(dmemXbar_io_in_2_req_ready),
    .io_in_2_req_valid(dmemXbar_io_in_2_req_valid),
    .io_in_2_req_bits_addr(dmemXbar_io_in_2_req_bits_addr),
    .io_in_2_req_bits_cmd(dmemXbar_io_in_2_req_bits_cmd),
    .io_in_2_req_bits_wdata(dmemXbar_io_in_2_req_bits_wdata),
    .io_in_2_resp_valid(dmemXbar_io_in_2_resp_valid),
    .io_in_2_resp_bits_rdata(dmemXbar_io_in_2_resp_bits_rdata),
    .io_out_req_ready(dmemXbar_io_out_req_ready),
    .io_out_req_valid(dmemXbar_io_out_req_valid),
    .io_out_req_bits_addr(dmemXbar_io_out_req_bits_addr),
    .io_out_req_bits_size(dmemXbar_io_out_req_bits_size),
    .io_out_req_bits_cmd(dmemXbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(dmemXbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(dmemXbar_io_out_req_bits_wdata),
    .io_out_resp_ready(dmemXbar_io_out_resp_ready),
    .io_out_resp_valid(dmemXbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(dmemXbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(dmemXbar_io_out_resp_bits_rdata)
  );
  EmbeddedTLB itlb ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
    .clock(itlb_clock),
    .reset(itlb_reset),
    .io_in_req_ready(itlb_io_in_req_ready),
    .io_in_req_valid(itlb_io_in_req_valid),
    .io_in_req_bits_addr(itlb_io_in_req_bits_addr),
    .io_in_req_bits_user(itlb_io_in_req_bits_user),
    .io_in_resp_ready(itlb_io_in_resp_ready),
    .io_in_resp_valid(itlb_io_in_resp_valid),
    .io_in_resp_bits_rdata(itlb_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(itlb_io_in_resp_bits_user),
    .io_out_req_ready(itlb_io_out_req_ready),
    .io_out_req_valid(itlb_io_out_req_valid),
    .io_out_req_bits_addr(itlb_io_out_req_bits_addr),
    .io_out_req_bits_user(itlb_io_out_req_bits_user),
    .io_out_resp_ready(itlb_io_out_resp_ready),
    .io_out_resp_valid(itlb_io_out_resp_valid),
    .io_out_resp_bits_rdata(itlb_io_out_resp_bits_rdata),
    .io_out_resp_bits_user(itlb_io_out_resp_bits_user),
    .io_mem_req_ready(itlb_io_mem_req_ready),
    .io_mem_req_valid(itlb_io_mem_req_valid),
    .io_mem_req_bits_addr(itlb_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(itlb_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(itlb_io_mem_req_bits_wdata),
    .io_mem_resp_valid(itlb_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(itlb_io_mem_resp_bits_rdata),
    .io_flush(itlb_io_flush),
    .io_csrMMU_priviledgeMode(itlb_io_csrMMU_priviledgeMode),
    .io_iaf(itlb_io_iaf),
    .CSRSATP(itlb_CSRSATP),
    .MOUFlushTLB(itlb_MOUFlushTLB)
  );
  PTERequestFilter filter ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
    .clock(filter_clock),
    .reset(filter_reset),
    .io_in_req_ready(filter_io_in_req_ready),
    .io_in_req_valid(filter_io_in_req_valid),
    .io_in_req_bits_addr(filter_io_in_req_bits_addr),
    .io_in_req_bits_cmd(filter_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(filter_io_in_req_bits_wdata),
    .io_in_resp_valid(filter_io_in_resp_valid),
    .io_in_resp_bits_rdata(filter_io_in_resp_bits_rdata),
    .io_out_req_ready(filter_io_out_req_ready),
    .io_out_req_valid(filter_io_out_req_valid),
    .io_out_req_bits_addr(filter_io_out_req_bits_addr),
    .io_out_req_bits_cmd(filter_io_out_req_bits_cmd),
    .io_out_req_bits_wdata(filter_io_out_req_bits_wdata),
    .io_out_resp_valid(filter_io_out_resp_valid),
    .io_out_resp_bits_rdata(filter_io_out_resp_bits_rdata),
    .io_u(filter_io_u)
  );
  Cache_fake io_imem_cache ( // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
    .clock(io_imem_cache_clock),
    .reset(io_imem_cache_reset),
    .io_in_req_ready(io_imem_cache_io_in_req_ready),
    .io_in_req_valid(io_imem_cache_io_in_req_valid),
    .io_in_req_bits_addr(io_imem_cache_io_in_req_bits_addr),
    .io_in_req_bits_user(io_imem_cache_io_in_req_bits_user),
    .io_in_resp_ready(io_imem_cache_io_in_resp_ready),
    .io_in_resp_valid(io_imem_cache_io_in_resp_valid),
    .io_in_resp_bits_rdata(io_imem_cache_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(io_imem_cache_io_in_resp_bits_user),
    .io_flush(io_imem_cache_io_flush),
    .io_out_mem_req_ready(io_imem_cache_io_out_mem_req_ready),
    .io_out_mem_req_valid(io_imem_cache_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(io_imem_cache_io_out_mem_req_bits_addr),
    .io_out_mem_resp_ready(io_imem_cache_io_out_mem_resp_ready),
    .io_out_mem_resp_valid(io_imem_cache_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_rdata(io_imem_cache_io_out_mem_resp_bits_rdata),
    .io_mmio_req_ready(io_imem_cache_io_mmio_req_ready),
    .io_mmio_req_valid(io_imem_cache_io_mmio_req_valid),
    .io_mmio_req_bits_addr(io_imem_cache_io_mmio_req_bits_addr),
    .io_mmio_resp_ready(io_imem_cache_io_mmio_resp_ready),
    .io_mmio_resp_valid(io_imem_cache_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(io_imem_cache_io_mmio_resp_bits_rdata)
  );
  EmbeddedTLB_1 dtlb ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 586:13]
    .clock(dtlb_clock),
    .reset(dtlb_reset),
    .io_in_req_ready(dtlb_io_in_req_ready),
    .io_in_req_valid(dtlb_io_in_req_valid),
    .io_in_req_bits_addr(dtlb_io_in_req_bits_addr),
    .io_in_req_bits_size(dtlb_io_in_req_bits_size),
    .io_in_req_bits_cmd(dtlb_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(dtlb_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(dtlb_io_in_req_bits_wdata),
    .io_in_resp_valid(dtlb_io_in_resp_valid),
    .io_in_resp_bits_rdata(dtlb_io_in_resp_bits_rdata),
    .io_out_req_ready(dtlb_io_out_req_ready),
    .io_out_req_valid(dtlb_io_out_req_valid),
    .io_out_req_bits_addr(dtlb_io_out_req_bits_addr),
    .io_out_req_bits_size(dtlb_io_out_req_bits_size),
    .io_out_req_bits_cmd(dtlb_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(dtlb_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(dtlb_io_out_req_bits_wdata),
    .io_out_resp_valid(dtlb_io_out_resp_valid),
    .io_out_resp_bits_rdata(dtlb_io_out_resp_bits_rdata),
    .io_mem_req_ready(dtlb_io_mem_req_ready),
    .io_mem_req_valid(dtlb_io_mem_req_valid),
    .io_mem_req_bits_addr(dtlb_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(dtlb_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(dtlb_io_mem_req_bits_wdata),
    .io_mem_resp_valid(dtlb_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(dtlb_io_mem_resp_bits_rdata),
    .io_csrMMU_priviledgeMode(dtlb_io_csrMMU_priviledgeMode),
    .io_csrMMU_status_sum(dtlb_io_csrMMU_status_sum),
    .io_csrMMU_status_mxr(dtlb_io_csrMMU_status_mxr),
    .io_csrMMU_loadPF(dtlb_io_csrMMU_loadPF),
    .io_csrMMU_storePF(dtlb_io_csrMMU_storePF),
    .io_csrMMU_laf(dtlb_io_csrMMU_laf),
    .io_csrMMU_saf(dtlb_io_csrMMU_saf),
    .lr(dtlb_lr),
    .scInflight(dtlb_scInflight),
    .amoReq(dtlb_amoReq),
    .lrAddr(dtlb_lrAddr),
    .paddr(dtlb_paddr),
    .CSRSATP(dtlb_CSRSATP),
    ._T_12_0(dtlb__T_12_0),
    .scIsSuccess_0(dtlb_scIsSuccess_0),
    .vmEnable_0(dtlb_vmEnable_0),
    .MOUFlushTLB(dtlb_MOUFlushTLB),
    .tlbFinish_0(dtlb_tlbFinish_0),
    ._T_13_1(dtlb__T_13_1)
  );
  PTERequestFilter_1 filter_1 ( // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 590:24]
    .clock(filter_1_clock),
    .reset(filter_1_reset),
    .io_in_req_ready(filter_1_io_in_req_ready),
    .io_in_req_valid(filter_1_io_in_req_valid),
    .io_in_req_bits_addr(filter_1_io_in_req_bits_addr),
    .io_in_req_bits_cmd(filter_1_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(filter_1_io_in_req_bits_wdata),
    .io_in_resp_valid(filter_1_io_in_resp_valid),
    .io_in_resp_bits_rdata(filter_1_io_in_resp_bits_rdata),
    .io_out_req_ready(filter_1_io_out_req_ready),
    .io_out_req_valid(filter_1_io_out_req_valid),
    .io_out_req_bits_addr(filter_1_io_out_req_bits_addr),
    .io_out_req_bits_cmd(filter_1_io_out_req_bits_cmd),
    .io_out_req_bits_wdata(filter_1_io_out_req_bits_wdata),
    .io_out_resp_valid(filter_1_io_out_resp_valid),
    .io_out_resp_bits_rdata(filter_1_io_out_resp_bits_rdata),
    .io_u(filter_1_io_u)
  );
  Cache_fake_1 io_dmem_cache ( // @[src/main/scala/nutcore/mem/Cache.scala 674:32]
    .clock(io_dmem_cache_clock),
    .reset(io_dmem_cache_reset),
    .io_in_req_ready(io_dmem_cache_io_in_req_ready),
    .io_in_req_valid(io_dmem_cache_io_in_req_valid),
    .io_in_req_bits_addr(io_dmem_cache_io_in_req_bits_addr),
    .io_in_req_bits_size(io_dmem_cache_io_in_req_bits_size),
    .io_in_req_bits_cmd(io_dmem_cache_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(io_dmem_cache_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(io_dmem_cache_io_in_req_bits_wdata),
    .io_in_resp_valid(io_dmem_cache_io_in_resp_valid),
    .io_in_resp_bits_cmd(io_dmem_cache_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(io_dmem_cache_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(io_dmem_cache_io_out_mem_req_ready),
    .io_out_mem_req_valid(io_dmem_cache_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(io_dmem_cache_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_size(io_dmem_cache_io_out_mem_req_bits_size),
    .io_out_mem_req_bits_cmd(io_dmem_cache_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wmask(io_dmem_cache_io_out_mem_req_bits_wmask),
    .io_out_mem_req_bits_wdata(io_dmem_cache_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_ready(io_dmem_cache_io_out_mem_resp_ready),
    .io_out_mem_resp_valid(io_dmem_cache_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(io_dmem_cache_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(io_dmem_cache_io_out_mem_resp_bits_rdata),
    .io_mmio_req_ready(io_dmem_cache_io_mmio_req_ready),
    .io_mmio_req_valid(io_dmem_cache_io_mmio_req_valid),
    .io_mmio_req_bits_addr(io_dmem_cache_io_mmio_req_bits_addr),
    .io_mmio_req_bits_cmd(io_dmem_cache_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(io_dmem_cache_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(io_dmem_cache_io_mmio_req_bits_wdata),
    .io_mmio_resp_ready(io_dmem_cache_io_mmio_resp_ready),
    .io_mmio_resp_valid(io_dmem_cache_io_mmio_resp_valid),
    .io_mmio_resp_bits_cmd(io_dmem_cache_io_mmio_resp_bits_cmd),
    .io_mmio_resp_bits_rdata(io_dmem_cache_io_mmio_resp_bits_rdata),
    .ismmio_0(io_dmem_cache_ismmio_0)
  );
  GEN_w64_toggle #(.COVER_INDEX(9135)) toggle_9135 (
    .clock(toggle_9135_clock),
    .reset(toggle_9135_reset),
    .valid(toggle_9135_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(9199)) toggle_9199 (
    .clock(toggle_9199_clock),
    .reset(toggle_9199_reset),
    .valid(toggle_9199_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(9238)) toggle_9238 (
    .clock(toggle_9238_clock),
    .reset(toggle_9238_reset),
    .valid(toggle_9238_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9277)) toggle_9277 (
    .clock(toggle_9277_clock),
    .reset(toggle_9277_reset),
    .valid(toggle_9277_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9278)) toggle_9278 (
    .clock(toggle_9278_clock),
    .reset(toggle_9278_reset),
    .valid(toggle_9278_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9279)) toggle_9279 (
    .clock(toggle_9279_clock),
    .reset(toggle_9279_reset),
    .valid(toggle_9279_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9280)) toggle_9280 (
    .clock(toggle_9280_clock),
    .reset(toggle_9280_reset),
    .valid(toggle_9280_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9281)) toggle_9281 (
    .clock(toggle_9281_clock),
    .reset(toggle_9281_reset),
    .valid(toggle_9281_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9282)) toggle_9282 (
    .clock(toggle_9282_clock),
    .reset(toggle_9282_reset),
    .valid(toggle_9282_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9283)) toggle_9283 (
    .clock(toggle_9283_clock),
    .reset(toggle_9283_reset),
    .valid(toggle_9283_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9284)) toggle_9284 (
    .clock(toggle_9284_clock),
    .reset(toggle_9284_reset),
    .valid(toggle_9284_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9285)) toggle_9285 (
    .clock(toggle_9285_clock),
    .reset(toggle_9285_reset),
    .valid(toggle_9285_valid)
  );
  GEN_w4_toggle #(.COVER_INDEX(9286)) toggle_9286 (
    .clock(toggle_9286_clock),
    .reset(toggle_9286_reset),
    .valid(toggle_9286_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9290)) toggle_9290 (
    .clock(toggle_9290_clock),
    .reset(toggle_9290_reset),
    .valid(toggle_9290_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9291)) toggle_9291 (
    .clock(toggle_9291_clock),
    .reset(toggle_9291_reset),
    .valid(toggle_9291_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9292)) toggle_9292 (
    .clock(toggle_9292_clock),
    .reset(toggle_9292_reset),
    .valid(toggle_9292_valid)
  );
  GEN_w3_toggle #(.COVER_INDEX(9293)) toggle_9293 (
    .clock(toggle_9293_clock),
    .reset(toggle_9293_reset),
    .valid(toggle_9293_valid)
  );
  GEN_w7_toggle #(.COVER_INDEX(9296)) toggle_9296 (
    .clock(toggle_9296_clock),
    .reset(toggle_9296_reset),
    .valid(toggle_9296_valid)
  );
  GEN_w5_toggle #(.COVER_INDEX(9303)) toggle_9303 (
    .clock(toggle_9303_clock),
    .reset(toggle_9303_reset),
    .valid(toggle_9303_valid)
  );
  GEN_w5_toggle #(.COVER_INDEX(9308)) toggle_9308 (
    .clock(toggle_9308_clock),
    .reset(toggle_9308_reset),
    .valid(toggle_9308_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9313)) toggle_9313 (
    .clock(toggle_9313_clock),
    .reset(toggle_9313_reset),
    .valid(toggle_9313_valid)
  );
  GEN_w5_toggle #(.COVER_INDEX(9314)) toggle_9314 (
    .clock(toggle_9314_clock),
    .reset(toggle_9314_reset),
    .valid(toggle_9314_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9319)) toggle_9319 (
    .clock(toggle_9319_clock),
    .reset(toggle_9319_reset),
    .valid(toggle_9319_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(9320)) toggle_9320 (
    .clock(toggle_9320_clock),
    .reset(toggle_9320_reset),
    .valid(toggle_9320_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(9384)) toggle_9384 (
    .clock(toggle_9384_clock),
    .reset(toggle_9384_reset),
    .valid(toggle_9384_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(9448)) toggle_9448 (
    .clock(toggle_9448_clock),
    .reset(toggle_9448_reset),
    .valid(toggle_9448_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(9487)) toggle_9487 (
    .clock(toggle_9487_clock),
    .reset(toggle_9487_reset),
    .valid(toggle_9487_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9526)) toggle_9526 (
    .clock(toggle_9526_clock),
    .reset(toggle_9526_reset),
    .valid(toggle_9526_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9527)) toggle_9527 (
    .clock(toggle_9527_clock),
    .reset(toggle_9527_reset),
    .valid(toggle_9527_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9528)) toggle_9528 (
    .clock(toggle_9528_clock),
    .reset(toggle_9528_reset),
    .valid(toggle_9528_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9529)) toggle_9529 (
    .clock(toggle_9529_clock),
    .reset(toggle_9529_reset),
    .valid(toggle_9529_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9530)) toggle_9530 (
    .clock(toggle_9530_clock),
    .reset(toggle_9530_reset),
    .valid(toggle_9530_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9531)) toggle_9531 (
    .clock(toggle_9531_clock),
    .reset(toggle_9531_reset),
    .valid(toggle_9531_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9532)) toggle_9532 (
    .clock(toggle_9532_clock),
    .reset(toggle_9532_reset),
    .valid(toggle_9532_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9533)) toggle_9533 (
    .clock(toggle_9533_clock),
    .reset(toggle_9533_reset),
    .valid(toggle_9533_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9534)) toggle_9534 (
    .clock(toggle_9534_clock),
    .reset(toggle_9534_reset),
    .valid(toggle_9534_valid)
  );
  GEN_w4_toggle #(.COVER_INDEX(9535)) toggle_9535 (
    .clock(toggle_9535_clock),
    .reset(toggle_9535_reset),
    .valid(toggle_9535_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9539)) toggle_9539 (
    .clock(toggle_9539_clock),
    .reset(toggle_9539_reset),
    .valid(toggle_9539_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9540)) toggle_9540 (
    .clock(toggle_9540_clock),
    .reset(toggle_9540_reset),
    .valid(toggle_9540_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9541)) toggle_9541 (
    .clock(toggle_9541_clock),
    .reset(toggle_9541_reset),
    .valid(toggle_9541_valid)
  );
  GEN_w3_toggle #(.COVER_INDEX(9542)) toggle_9542 (
    .clock(toggle_9542_clock),
    .reset(toggle_9542_reset),
    .valid(toggle_9542_valid)
  );
  GEN_w7_toggle #(.COVER_INDEX(9545)) toggle_9545 (
    .clock(toggle_9545_clock),
    .reset(toggle_9545_reset),
    .valid(toggle_9545_valid)
  );
  GEN_w5_toggle #(.COVER_INDEX(9552)) toggle_9552 (
    .clock(toggle_9552_clock),
    .reset(toggle_9552_reset),
    .valid(toggle_9552_valid)
  );
  GEN_w5_toggle #(.COVER_INDEX(9557)) toggle_9557 (
    .clock(toggle_9557_clock),
    .reset(toggle_9557_reset),
    .valid(toggle_9557_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9562)) toggle_9562 (
    .clock(toggle_9562_clock),
    .reset(toggle_9562_reset),
    .valid(toggle_9562_valid)
  );
  GEN_w5_toggle #(.COVER_INDEX(9563)) toggle_9563 (
    .clock(toggle_9563_clock),
    .reset(toggle_9563_reset),
    .valid(toggle_9563_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9568)) toggle_9568 (
    .clock(toggle_9568_clock),
    .reset(toggle_9568_reset),
    .valid(toggle_9568_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(9569)) toggle_9569 (
    .clock(toggle_9569_clock),
    .reset(toggle_9569_reset),
    .valid(toggle_9569_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(9633)) toggle_9633 (
    .clock(toggle_9633_clock),
    .reset(toggle_9633_reset),
    .valid(toggle_9633_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(9697)) toggle_9697 (
    .clock(toggle_9697_clock),
    .reset(toggle_9697_reset),
    .valid(toggle_9697_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(9736)) toggle_9736 (
    .clock(toggle_9736_clock),
    .reset(toggle_9736_reset),
    .valid(toggle_9736_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9775)) toggle_9775 (
    .clock(toggle_9775_clock),
    .reset(toggle_9775_reset),
    .valid(toggle_9775_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9776)) toggle_9776 (
    .clock(toggle_9776_clock),
    .reset(toggle_9776_reset),
    .valid(toggle_9776_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9777)) toggle_9777 (
    .clock(toggle_9777_clock),
    .reset(toggle_9777_reset),
    .valid(toggle_9777_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9778)) toggle_9778 (
    .clock(toggle_9778_clock),
    .reset(toggle_9778_reset),
    .valid(toggle_9778_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9779)) toggle_9779 (
    .clock(toggle_9779_clock),
    .reset(toggle_9779_reset),
    .valid(toggle_9779_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9780)) toggle_9780 (
    .clock(toggle_9780_clock),
    .reset(toggle_9780_reset),
    .valid(toggle_9780_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9781)) toggle_9781 (
    .clock(toggle_9781_clock),
    .reset(toggle_9781_reset),
    .valid(toggle_9781_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9782)) toggle_9782 (
    .clock(toggle_9782_clock),
    .reset(toggle_9782_reset),
    .valid(toggle_9782_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9783)) toggle_9783 (
    .clock(toggle_9783_clock),
    .reset(toggle_9783_reset),
    .valid(toggle_9783_valid)
  );
  GEN_w4_toggle #(.COVER_INDEX(9784)) toggle_9784 (
    .clock(toggle_9784_clock),
    .reset(toggle_9784_reset),
    .valid(toggle_9784_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9788)) toggle_9788 (
    .clock(toggle_9788_clock),
    .reset(toggle_9788_reset),
    .valid(toggle_9788_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9789)) toggle_9789 (
    .clock(toggle_9789_clock),
    .reset(toggle_9789_reset),
    .valid(toggle_9789_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9790)) toggle_9790 (
    .clock(toggle_9790_clock),
    .reset(toggle_9790_reset),
    .valid(toggle_9790_valid)
  );
  GEN_w3_toggle #(.COVER_INDEX(9791)) toggle_9791 (
    .clock(toggle_9791_clock),
    .reset(toggle_9791_reset),
    .valid(toggle_9791_valid)
  );
  GEN_w7_toggle #(.COVER_INDEX(9794)) toggle_9794 (
    .clock(toggle_9794_clock),
    .reset(toggle_9794_reset),
    .valid(toggle_9794_valid)
  );
  GEN_w5_toggle #(.COVER_INDEX(9801)) toggle_9801 (
    .clock(toggle_9801_clock),
    .reset(toggle_9801_reset),
    .valid(toggle_9801_valid)
  );
  GEN_w5_toggle #(.COVER_INDEX(9806)) toggle_9806 (
    .clock(toggle_9806_clock),
    .reset(toggle_9806_reset),
    .valid(toggle_9806_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9811)) toggle_9811 (
    .clock(toggle_9811_clock),
    .reset(toggle_9811_reset),
    .valid(toggle_9811_valid)
  );
  GEN_w5_toggle #(.COVER_INDEX(9812)) toggle_9812 (
    .clock(toggle_9812_clock),
    .reset(toggle_9812_reset),
    .valid(toggle_9812_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(9817)) toggle_9817 (
    .clock(toggle_9817_clock),
    .reset(toggle_9817_reset),
    .valid(toggle_9817_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(9818)) toggle_9818 (
    .clock(toggle_9818_clock),
    .reset(toggle_9818_reset),
    .valid(toggle_9818_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(9882)) toggle_9882 (
    .clock(toggle_9882_clock),
    .reset(toggle_9882_reset),
    .valid(toggle_9882_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(9946)) toggle_9946 (
    .clock(toggle_9946_clock),
    .reset(toggle_9946_reset),
    .valid(toggle_9946_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(9985)) toggle_9985 (
    .clock(toggle_9985_clock),
    .reset(toggle_9985_reset),
    .valid(toggle_9985_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10024)) toggle_10024 (
    .clock(toggle_10024_clock),
    .reset(toggle_10024_reset),
    .valid(toggle_10024_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10025)) toggle_10025 (
    .clock(toggle_10025_clock),
    .reset(toggle_10025_reset),
    .valid(toggle_10025_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10026)) toggle_10026 (
    .clock(toggle_10026_clock),
    .reset(toggle_10026_reset),
    .valid(toggle_10026_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10027)) toggle_10027 (
    .clock(toggle_10027_clock),
    .reset(toggle_10027_reset),
    .valid(toggle_10027_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10028)) toggle_10028 (
    .clock(toggle_10028_clock),
    .reset(toggle_10028_reset),
    .valid(toggle_10028_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10029)) toggle_10029 (
    .clock(toggle_10029_clock),
    .reset(toggle_10029_reset),
    .valid(toggle_10029_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10030)) toggle_10030 (
    .clock(toggle_10030_clock),
    .reset(toggle_10030_reset),
    .valid(toggle_10030_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10031)) toggle_10031 (
    .clock(toggle_10031_clock),
    .reset(toggle_10031_reset),
    .valid(toggle_10031_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10032)) toggle_10032 (
    .clock(toggle_10032_clock),
    .reset(toggle_10032_reset),
    .valid(toggle_10032_valid)
  );
  GEN_w4_toggle #(.COVER_INDEX(10033)) toggle_10033 (
    .clock(toggle_10033_clock),
    .reset(toggle_10033_reset),
    .valid(toggle_10033_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10037)) toggle_10037 (
    .clock(toggle_10037_clock),
    .reset(toggle_10037_reset),
    .valid(toggle_10037_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10038)) toggle_10038 (
    .clock(toggle_10038_clock),
    .reset(toggle_10038_reset),
    .valid(toggle_10038_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10039)) toggle_10039 (
    .clock(toggle_10039_clock),
    .reset(toggle_10039_reset),
    .valid(toggle_10039_valid)
  );
  GEN_w3_toggle #(.COVER_INDEX(10040)) toggle_10040 (
    .clock(toggle_10040_clock),
    .reset(toggle_10040_reset),
    .valid(toggle_10040_valid)
  );
  GEN_w7_toggle #(.COVER_INDEX(10043)) toggle_10043 (
    .clock(toggle_10043_clock),
    .reset(toggle_10043_reset),
    .valid(toggle_10043_valid)
  );
  GEN_w5_toggle #(.COVER_INDEX(10050)) toggle_10050 (
    .clock(toggle_10050_clock),
    .reset(toggle_10050_reset),
    .valid(toggle_10050_valid)
  );
  GEN_w5_toggle #(.COVER_INDEX(10055)) toggle_10055 (
    .clock(toggle_10055_clock),
    .reset(toggle_10055_reset),
    .valid(toggle_10055_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10060)) toggle_10060 (
    .clock(toggle_10060_clock),
    .reset(toggle_10060_reset),
    .valid(toggle_10060_valid)
  );
  GEN_w5_toggle #(.COVER_INDEX(10061)) toggle_10061 (
    .clock(toggle_10061_clock),
    .reset(toggle_10061_reset),
    .valid(toggle_10061_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10066)) toggle_10066 (
    .clock(toggle_10066_clock),
    .reset(toggle_10066_reset),
    .valid(toggle_10066_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(10067)) toggle_10067 (
    .clock(toggle_10067_clock),
    .reset(toggle_10067_reset),
    .valid(toggle_10067_valid)
  );
  GEN_w2_toggle #(.COVER_INDEX(10131)) toggle_10131 (
    .clock(toggle_10131_clock),
    .reset(toggle_10131_reset),
    .valid(toggle_10131_valid)
  );
  GEN_w2_toggle #(.COVER_INDEX(10133)) toggle_10133 (
    .clock(toggle_10133_clock),
    .reset(toggle_10133_reset),
    .valid(toggle_10133_valid)
  );
  assign io_imem_mem_req_valid = io_imem_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/NutCore.scala 190:13]
  assign io_imem_mem_req_bits_addr = io_imem_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 190:13]
  assign io_dmem_mem_req_valid = io_dmem_cache_io_out_mem_req_valid; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_mem_req_bits_addr = io_dmem_cache_io_out_mem_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_mem_req_bits_size = io_dmem_cache_io_out_mem_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_mem_req_bits_cmd = io_dmem_cache_io_out_mem_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_mem_req_bits_wmask = io_dmem_cache_io_out_mem_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_mem_req_bits_wdata = io_dmem_cache_io_out_mem_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_mmio_req_valid = mmioXbar_io_out_req_valid; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign io_mmio_req_bits_addr = mmioXbar_io_out_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign io_mmio_req_bits_cmd = mmioXbar_io_out_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign io_mmio_req_bits_wmask = mmioXbar_io_out_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign io_mmio_req_bits_wdata = mmioXbar_io_out_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign isWFI = frontend_isWFI;
  assign frontend_clock = clock;
  assign frontend_reset = reset;
  assign frontend_io_imem_req_ready = itlb_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign frontend_io_imem_resp_valid = itlb_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign frontend_io_imem_resp_bits_rdata = itlb_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign frontend_io_imem_resp_bits_user = itlb_io_in_resp_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign frontend_io_out_0_ready = ringBufferAllowin | ~frontend_io_out_0_valid; // @[src/main/scala/utils/PipelineVector.scala 50:36]
  assign frontend_io_redirect_target = backend_io_redirect_target; // @[src/main/scala/nutcore/NutCore.scala 218:26]
  assign frontend_io_redirect_valid = backend_io_redirect_valid; // @[src/main/scala/nutcore/NutCore.scala 218:26]
  assign frontend_io_iaf = itlb_io_iaf; // @[src/main/scala/nutcore/NutCore.scala 189:21]
  assign frontend_io_sfence_vma_invalid = backend_io_sfence_vma_invalid; // @[src/main/scala/nutcore/NutCore.scala 215:36]
  assign frontend_io_wfi_invalid = backend_io_wfi_invalid; // @[src/main/scala/nutcore/NutCore.scala 216:29]
  assign frontend_REG_valid = backend_REG_valid;
  assign frontend_REG_pc = backend_REG_pc;
  assign frontend_REG_isMissPredict = backend_REG_isMissPredict;
  assign frontend_REG_actualTarget = backend_REG_actualTarget;
  assign frontend_REG_fuOpType = backend_REG_fuOpType;
  assign frontend_REG_btbType = backend_REG_btbType;
  assign frontend_REG_isRVC = backend_REG_isRVC;
  assign frontend_flushICache = backend_flushICache;
  assign frontend_flushTLB = backend_flushTLB;
  assign frontend_intrVecIDU = backend_intrVecIDU;
  assign backend_clock = clock;
  assign backend_reset = reset;
  assign backend_io_in_0_valid = ringBufferHead != ringBufferTail; // @[src/main/scala/utils/PipelineVector.scala 56:34]
  assign backend_io_in_0_bits_cf_instr = 2'h3 == ringBufferTail ? dataBuffer_3_cf_instr : _GEN_1343; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_pc = 2'h3 == ringBufferTail ? dataBuffer_3_cf_pc : _GEN_1339; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_pnpc = 2'h3 == ringBufferTail ? dataBuffer_3_cf_pnpc : _GEN_1335; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_exceptionVec_1 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_exceptionVec_1 : _GEN_1263; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_exceptionVec_2 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_exceptionVec_2 : _GEN_1267; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_exceptionVec_12 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_exceptionVec_12 : _GEN_1307; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_1 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_1 : _GEN_1215; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_3 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_3 : _GEN_1223; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_5 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_5 : _GEN_1231; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_7 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_7 : _GEN_1239; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_9 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_9 : _GEN_1247; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_intrVec_11 = 2'h3 == ringBufferTail ? dataBuffer_3_cf_intrVec_11 : _GEN_1255; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_brIdx = 2'h3 == ringBufferTail ? dataBuffer_3_cf_brIdx : _GEN_1207; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_cf_crossBoundaryFault = 2'h3 == ringBufferTail ? dataBuffer_3_cf_crossBoundaryFault :
    _GEN_1199; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_src1Type = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_src1Type : _GEN_1183; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_src2Type = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_src2Type : _GEN_1179; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_fuType = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_fuType : _GEN_1175; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_fuOpType = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_fuOpType : _GEN_1171; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfSrc1 = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_rfSrc1 : _GEN_1167; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfSrc2 = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_rfSrc2 : _GEN_1163; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfWen = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_rfWen : _GEN_1159; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_rfDest = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_rfDest : _GEN_1155; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_ctrl_isNutCoreTrap = 2'h3 == ringBufferTail ? dataBuffer_3_ctrl_isNutCoreTrap : _GEN_1151; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_in_0_bits_data_imm = 2'h3 == ringBufferTail ? dataBuffer_3_data_imm : _GEN_1123; // @[src/main/scala/utils/PipelineVector.scala 55:{15,15}]
  assign backend_io_flush = frontend_io_flushVec[3:2]; // @[src/main/scala/nutcore/NutCore.scala 219:45]
  assign backend_io_dmem_req_ready = dtlb_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign backend_io_dmem_resp_valid = dtlb_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign backend_io_dmem_resp_bits_rdata = dtlb_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign backend_io_memMMU_dmem_loadPF = dtlb_io_csrMMU_loadPF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign backend_io_memMMU_dmem_storePF = dtlb_io_csrMMU_storePF; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign backend_io_memMMU_dmem_laf = dtlb_io_csrMMU_laf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign backend_io_memMMU_dmem_saf = dtlb_io_csrMMU_saf; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign backend_io_extra_meip_0 = io_extra_meip_0;
  assign backend_paddr = dtlb_paddr;
  assign backend__T_12 = dtlb__T_12_0;
  assign backend_scIsSuccess = dtlb_scIsSuccess_0;
  assign backend_io_extra_mtip = io_extra_mtip;
  assign backend_vmEnable = dtlb_vmEnable_0;
  assign backend_tlbFinish = dtlb_tlbFinish_0;
  assign backend_ismmio = io_dmem_cache_ismmio_0;
  assign backend__T_13_0 = dtlb__T_13_1;
  assign backend_io_extra_msip = io_extra_msip;
  assign mmioXbar_clock = clock;
  assign mmioXbar_reset = reset;
  assign mmioXbar_io_in_0_req_valid = io_imem_cache_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_0_req_bits_addr = io_imem_cache_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_valid = io_dmem_cache_io_mmio_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_bits_addr = io_dmem_cache_io_mmio_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_bits_cmd = io_dmem_cache_io_mmio_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_bits_wmask = io_dmem_cache_io_mmio_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_in_1_req_bits_wdata = io_dmem_cache_io_mmio_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign mmioXbar_io_out_req_ready = io_mmio_req_ready; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign mmioXbar_io_out_resp_valid = io_mmio_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign mmioXbar_io_out_resp_bits_cmd = io_mmio_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign mmioXbar_io_out_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 224:13]
  assign dmemXbar_clock = clock;
  assign dmemXbar_reset = reset;
  assign dmemXbar_io_in_0_req_valid = dtlb_io_out_req_valid; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_0_req_bits_addr = dtlb_io_out_req_bits_addr; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_0_req_bits_size = dtlb_io_out_req_bits_size; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_0_req_bits_cmd = dtlb_io_out_req_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_0_req_bits_wmask = dtlb_io_out_req_bits_wmask; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_0_req_bits_wdata = dtlb_io_out_req_bits_wdata; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dmemXbar_io_in_1_req_valid = filter_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_1_req_bits_addr = filter_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_1_req_bits_cmd = filter_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_1_req_bits_wdata = filter_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_2_req_valid = filter_1_io_out_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_2_req_bits_addr = filter_1_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_2_req_bits_cmd = filter_1_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_in_2_req_bits_wdata = filter_1_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign dmemXbar_io_out_req_ready = io_dmem_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign dmemXbar_io_out_resp_valid = io_dmem_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign dmemXbar_io_out_resp_bits_cmd = io_dmem_cache_io_in_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign dmemXbar_io_out_resp_bits_rdata = io_dmem_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign itlb_clock = clock;
  assign itlb_reset = reset;
  assign itlb_io_in_req_valid = frontend_io_imem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign itlb_io_in_req_bits_addr = frontend_io_imem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign itlb_io_in_req_bits_user = frontend_io_imem_req_bits_user; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign itlb_io_in_resp_ready = frontend_io_imem_resp_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign itlb_io_out_req_ready = io_imem_cache_io_in_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign itlb_io_out_resp_valid = io_imem_cache_io_in_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign itlb_io_out_resp_bits_rdata = io_imem_cache_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign itlb_io_out_resp_bits_user = io_imem_cache_io_in_resp_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign itlb_io_mem_req_ready = filter_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign itlb_io_mem_resp_valid = filter_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign itlb_io_mem_resp_bits_rdata = filter_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign itlb_io_flush = frontend_io_flushVec[0]; // @[src/main/scala/nutcore/NutCore.scala 184:35]
  assign itlb_io_csrMMU_priviledgeMode = backend_io_memMMU_imem_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign itlb_CSRSATP = backend_satp;
  assign itlb_MOUFlushTLB = backend_flushTLB;
  assign filter_clock = clock;
  assign filter_reset = reset;
  assign filter_io_in_req_valid = itlb_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_io_in_req_bits_addr = itlb_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_io_in_req_bits_cmd = itlb_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_io_in_req_bits_wdata = itlb_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_io_out_req_ready = dmemXbar_io_in_1_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign filter_io_out_resp_valid = dmemXbar_io_in_1_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign filter_io_out_resp_bits_rdata = dmemXbar_io_in_1_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign filter_io_u = backend_io_memMMU_imem_priviledgeMode == 2'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 591:42]
  assign io_imem_cache_clock = clock;
  assign io_imem_cache_reset = reset;
  assign io_imem_cache_io_in_req_valid = itlb_io_out_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_imem_cache_io_in_req_bits_addr = itlb_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_imem_cache_io_in_req_bits_user = itlb_io_out_req_bits_user; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_imem_cache_io_in_resp_ready = itlb_io_out_resp_ready; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_imem_cache_io_flush = frontend_io_flushVec[0] ? 2'h3 : 2'h0; // @[src/main/scala/nutcore/NutCore.scala 193:19]
  assign io_imem_cache_io_out_mem_req_ready = io_imem_mem_req_ready; // @[src/main/scala/nutcore/NutCore.scala 190:13]
  assign io_imem_cache_io_out_mem_resp_valid = io_imem_mem_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 190:13]
  assign io_imem_cache_io_out_mem_resp_bits_rdata = io_imem_mem_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 190:13]
  assign io_imem_cache_io_mmio_req_ready = mmioXbar_io_in_0_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign io_imem_cache_io_mmio_resp_valid = mmioXbar_io_in_0_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign io_imem_cache_io_mmio_resp_bits_rdata = mmioXbar_io_in_0_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign dtlb_clock = clock;
  assign dtlb_reset = reset;
  assign dtlb_io_in_req_valid = backend_io_dmem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign dtlb_io_in_req_bits_addr = backend_io_dmem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign dtlb_io_in_req_bits_size = backend_io_dmem_req_bits_size; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign dtlb_io_in_req_bits_cmd = backend_io_dmem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign dtlb_io_in_req_bits_wmask = backend_io_dmem_req_bits_wmask; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign dtlb_io_in_req_bits_wdata = backend_io_dmem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 592:15]
  assign dtlb_io_out_req_ready = dmemXbar_io_in_0_req_ready; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dtlb_io_out_resp_valid = dmemXbar_io_in_0_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dtlb_io_out_resp_bits_rdata = dmemXbar_io_in_0_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 206:23]
  assign dtlb_io_mem_req_ready = filter_1_io_in_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign dtlb_io_mem_resp_valid = filter_1_io_in_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign dtlb_io_mem_resp_bits_rdata = filter_1_io_in_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign dtlb_io_csrMMU_priviledgeMode = backend_io_memMMU_dmem_priviledgeMode; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign dtlb_io_csrMMU_status_sum = backend_io_memMMU_dmem_status_sum; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign dtlb_io_csrMMU_status_mxr = backend_io_memMMU_dmem_status_mxr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 596:19]
  assign dtlb_lr = backend_lr;
  assign dtlb_scInflight = backend_scInflight;
  assign dtlb_amoReq = backend_amoReq;
  assign dtlb_lrAddr = backend_lrAddr;
  assign dtlb_CSRSATP = backend_satp;
  assign dtlb_MOUFlushTLB = backend_flushTLB;
  assign filter_1_clock = clock;
  assign filter_1_reset = reset;
  assign filter_1_io_in_req_valid = dtlb_io_mem_req_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_1_io_in_req_bits_addr = dtlb_io_mem_req_bits_addr; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_1_io_in_req_bits_cmd = dtlb_io_mem_req_bits_cmd; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_1_io_in_req_bits_wdata = dtlb_io_mem_req_bits_wdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 593:16]
  assign filter_1_io_out_req_ready = dmemXbar_io_in_2_req_ready; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign filter_1_io_out_resp_valid = dmemXbar_io_in_2_resp_valid; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign filter_1_io_out_resp_bits_rdata = dmemXbar_io_in_2_resp_bits_rdata; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 594:19]
  assign filter_1_io_u = backend_io_memMMU_dmem_priviledgeMode == 2'h0; // @[src/main/scala/nutcore/mem/EmbeddedTLB.scala 591:42]
  assign io_dmem_cache_clock = clock;
  assign io_dmem_cache_reset = reset;
  assign io_dmem_cache_io_in_req_valid = dmemXbar_io_out_req_valid; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_req_bits_addr = dmemXbar_io_out_req_bits_addr; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_req_bits_size = dmemXbar_io_out_req_bits_size; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_req_bits_cmd = dmemXbar_io_out_req_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_req_bits_wmask = dmemXbar_io_out_req_bits_wmask; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_in_req_bits_wdata = dmemXbar_io_out_req_bits_wdata; // @[src/main/scala/nutcore/mem/Cache.scala 676:17]
  assign io_dmem_cache_io_out_mem_req_ready = io_dmem_mem_req_ready; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_cache_io_out_mem_resp_valid = io_dmem_mem_resp_valid; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_cache_io_out_mem_resp_bits_cmd = io_dmem_mem_resp_bits_cmd; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_cache_io_out_mem_resp_bits_rdata = io_dmem_mem_resp_bits_rdata; // @[src/main/scala/nutcore/NutCore.scala 207:13]
  assign io_dmem_cache_io_mmio_req_ready = mmioXbar_io_in_1_req_ready; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign io_dmem_cache_io_mmio_resp_valid = mmioXbar_io_in_1_resp_valid; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign io_dmem_cache_io_mmio_resp_bits_cmd = mmioXbar_io_in_1_resp_bits_cmd; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign io_dmem_cache_io_mmio_resp_bits_rdata = mmioXbar_io_in_1_resp_bits_rdata; // @[src/main/scala/nutcore/mem/Cache.scala 677:13]
  assign toggle_9135_clock = clock;
  assign toggle_9135_reset = reset;
  assign toggle_9135_valid = dataBuffer_0_cf_instr ^ toggle_9135_valid_reg;
  assign toggle_9199_clock = clock;
  assign toggle_9199_reset = reset;
  assign toggle_9199_valid = dataBuffer_0_cf_pc ^ toggle_9199_valid_reg;
  assign toggle_9238_clock = clock;
  assign toggle_9238_reset = reset;
  assign toggle_9238_valid = dataBuffer_0_cf_pnpc ^ toggle_9238_valid_reg;
  assign toggle_9277_clock = clock;
  assign toggle_9277_reset = reset;
  assign toggle_9277_valid = dataBuffer_0_cf_exceptionVec_1 ^ toggle_9277_valid_reg;
  assign toggle_9278_clock = clock;
  assign toggle_9278_reset = reset;
  assign toggle_9278_valid = dataBuffer_0_cf_exceptionVec_2 ^ toggle_9278_valid_reg;
  assign toggle_9279_clock = clock;
  assign toggle_9279_reset = reset;
  assign toggle_9279_valid = dataBuffer_0_cf_exceptionVec_12 ^ toggle_9279_valid_reg;
  assign toggle_9280_clock = clock;
  assign toggle_9280_reset = reset;
  assign toggle_9280_valid = dataBuffer_0_cf_intrVec_1 ^ toggle_9280_valid_reg;
  assign toggle_9281_clock = clock;
  assign toggle_9281_reset = reset;
  assign toggle_9281_valid = dataBuffer_0_cf_intrVec_3 ^ toggle_9281_valid_reg;
  assign toggle_9282_clock = clock;
  assign toggle_9282_reset = reset;
  assign toggle_9282_valid = dataBuffer_0_cf_intrVec_5 ^ toggle_9282_valid_reg;
  assign toggle_9283_clock = clock;
  assign toggle_9283_reset = reset;
  assign toggle_9283_valid = dataBuffer_0_cf_intrVec_7 ^ toggle_9283_valid_reg;
  assign toggle_9284_clock = clock;
  assign toggle_9284_reset = reset;
  assign toggle_9284_valid = dataBuffer_0_cf_intrVec_9 ^ toggle_9284_valid_reg;
  assign toggle_9285_clock = clock;
  assign toggle_9285_reset = reset;
  assign toggle_9285_valid = dataBuffer_0_cf_intrVec_11 ^ toggle_9285_valid_reg;
  assign toggle_9286_clock = clock;
  assign toggle_9286_reset = reset;
  assign toggle_9286_valid = dataBuffer_0_cf_brIdx ^ toggle_9286_valid_reg;
  assign toggle_9290_clock = clock;
  assign toggle_9290_reset = reset;
  assign toggle_9290_valid = dataBuffer_0_cf_crossBoundaryFault ^ toggle_9290_valid_reg;
  assign toggle_9291_clock = clock;
  assign toggle_9291_reset = reset;
  assign toggle_9291_valid = dataBuffer_0_ctrl_src1Type ^ toggle_9291_valid_reg;
  assign toggle_9292_clock = clock;
  assign toggle_9292_reset = reset;
  assign toggle_9292_valid = dataBuffer_0_ctrl_src2Type ^ toggle_9292_valid_reg;
  assign toggle_9293_clock = clock;
  assign toggle_9293_reset = reset;
  assign toggle_9293_valid = dataBuffer_0_ctrl_fuType ^ toggle_9293_valid_reg;
  assign toggle_9296_clock = clock;
  assign toggle_9296_reset = reset;
  assign toggle_9296_valid = dataBuffer_0_ctrl_fuOpType ^ toggle_9296_valid_reg;
  assign toggle_9303_clock = clock;
  assign toggle_9303_reset = reset;
  assign toggle_9303_valid = dataBuffer_0_ctrl_rfSrc1 ^ toggle_9303_valid_reg;
  assign toggle_9308_clock = clock;
  assign toggle_9308_reset = reset;
  assign toggle_9308_valid = dataBuffer_0_ctrl_rfSrc2 ^ toggle_9308_valid_reg;
  assign toggle_9313_clock = clock;
  assign toggle_9313_reset = reset;
  assign toggle_9313_valid = dataBuffer_0_ctrl_rfWen ^ toggle_9313_valid_reg;
  assign toggle_9314_clock = clock;
  assign toggle_9314_reset = reset;
  assign toggle_9314_valid = dataBuffer_0_ctrl_rfDest ^ toggle_9314_valid_reg;
  assign toggle_9319_clock = clock;
  assign toggle_9319_reset = reset;
  assign toggle_9319_valid = dataBuffer_0_ctrl_isNutCoreTrap ^ toggle_9319_valid_reg;
  assign toggle_9320_clock = clock;
  assign toggle_9320_reset = reset;
  assign toggle_9320_valid = dataBuffer_0_data_imm ^ toggle_9320_valid_reg;
  assign toggle_9384_clock = clock;
  assign toggle_9384_reset = reset;
  assign toggle_9384_valid = dataBuffer_1_cf_instr ^ toggle_9384_valid_reg;
  assign toggle_9448_clock = clock;
  assign toggle_9448_reset = reset;
  assign toggle_9448_valid = dataBuffer_1_cf_pc ^ toggle_9448_valid_reg;
  assign toggle_9487_clock = clock;
  assign toggle_9487_reset = reset;
  assign toggle_9487_valid = dataBuffer_1_cf_pnpc ^ toggle_9487_valid_reg;
  assign toggle_9526_clock = clock;
  assign toggle_9526_reset = reset;
  assign toggle_9526_valid = dataBuffer_1_cf_exceptionVec_1 ^ toggle_9526_valid_reg;
  assign toggle_9527_clock = clock;
  assign toggle_9527_reset = reset;
  assign toggle_9527_valid = dataBuffer_1_cf_exceptionVec_2 ^ toggle_9527_valid_reg;
  assign toggle_9528_clock = clock;
  assign toggle_9528_reset = reset;
  assign toggle_9528_valid = dataBuffer_1_cf_exceptionVec_12 ^ toggle_9528_valid_reg;
  assign toggle_9529_clock = clock;
  assign toggle_9529_reset = reset;
  assign toggle_9529_valid = dataBuffer_1_cf_intrVec_1 ^ toggle_9529_valid_reg;
  assign toggle_9530_clock = clock;
  assign toggle_9530_reset = reset;
  assign toggle_9530_valid = dataBuffer_1_cf_intrVec_3 ^ toggle_9530_valid_reg;
  assign toggle_9531_clock = clock;
  assign toggle_9531_reset = reset;
  assign toggle_9531_valid = dataBuffer_1_cf_intrVec_5 ^ toggle_9531_valid_reg;
  assign toggle_9532_clock = clock;
  assign toggle_9532_reset = reset;
  assign toggle_9532_valid = dataBuffer_1_cf_intrVec_7 ^ toggle_9532_valid_reg;
  assign toggle_9533_clock = clock;
  assign toggle_9533_reset = reset;
  assign toggle_9533_valid = dataBuffer_1_cf_intrVec_9 ^ toggle_9533_valid_reg;
  assign toggle_9534_clock = clock;
  assign toggle_9534_reset = reset;
  assign toggle_9534_valid = dataBuffer_1_cf_intrVec_11 ^ toggle_9534_valid_reg;
  assign toggle_9535_clock = clock;
  assign toggle_9535_reset = reset;
  assign toggle_9535_valid = dataBuffer_1_cf_brIdx ^ toggle_9535_valid_reg;
  assign toggle_9539_clock = clock;
  assign toggle_9539_reset = reset;
  assign toggle_9539_valid = dataBuffer_1_cf_crossBoundaryFault ^ toggle_9539_valid_reg;
  assign toggle_9540_clock = clock;
  assign toggle_9540_reset = reset;
  assign toggle_9540_valid = dataBuffer_1_ctrl_src1Type ^ toggle_9540_valid_reg;
  assign toggle_9541_clock = clock;
  assign toggle_9541_reset = reset;
  assign toggle_9541_valid = dataBuffer_1_ctrl_src2Type ^ toggle_9541_valid_reg;
  assign toggle_9542_clock = clock;
  assign toggle_9542_reset = reset;
  assign toggle_9542_valid = dataBuffer_1_ctrl_fuType ^ toggle_9542_valid_reg;
  assign toggle_9545_clock = clock;
  assign toggle_9545_reset = reset;
  assign toggle_9545_valid = dataBuffer_1_ctrl_fuOpType ^ toggle_9545_valid_reg;
  assign toggle_9552_clock = clock;
  assign toggle_9552_reset = reset;
  assign toggle_9552_valid = dataBuffer_1_ctrl_rfSrc1 ^ toggle_9552_valid_reg;
  assign toggle_9557_clock = clock;
  assign toggle_9557_reset = reset;
  assign toggle_9557_valid = dataBuffer_1_ctrl_rfSrc2 ^ toggle_9557_valid_reg;
  assign toggle_9562_clock = clock;
  assign toggle_9562_reset = reset;
  assign toggle_9562_valid = dataBuffer_1_ctrl_rfWen ^ toggle_9562_valid_reg;
  assign toggle_9563_clock = clock;
  assign toggle_9563_reset = reset;
  assign toggle_9563_valid = dataBuffer_1_ctrl_rfDest ^ toggle_9563_valid_reg;
  assign toggle_9568_clock = clock;
  assign toggle_9568_reset = reset;
  assign toggle_9568_valid = dataBuffer_1_ctrl_isNutCoreTrap ^ toggle_9568_valid_reg;
  assign toggle_9569_clock = clock;
  assign toggle_9569_reset = reset;
  assign toggle_9569_valid = dataBuffer_1_data_imm ^ toggle_9569_valid_reg;
  assign toggle_9633_clock = clock;
  assign toggle_9633_reset = reset;
  assign toggle_9633_valid = dataBuffer_2_cf_instr ^ toggle_9633_valid_reg;
  assign toggle_9697_clock = clock;
  assign toggle_9697_reset = reset;
  assign toggle_9697_valid = dataBuffer_2_cf_pc ^ toggle_9697_valid_reg;
  assign toggle_9736_clock = clock;
  assign toggle_9736_reset = reset;
  assign toggle_9736_valid = dataBuffer_2_cf_pnpc ^ toggle_9736_valid_reg;
  assign toggle_9775_clock = clock;
  assign toggle_9775_reset = reset;
  assign toggle_9775_valid = dataBuffer_2_cf_exceptionVec_1 ^ toggle_9775_valid_reg;
  assign toggle_9776_clock = clock;
  assign toggle_9776_reset = reset;
  assign toggle_9776_valid = dataBuffer_2_cf_exceptionVec_2 ^ toggle_9776_valid_reg;
  assign toggle_9777_clock = clock;
  assign toggle_9777_reset = reset;
  assign toggle_9777_valid = dataBuffer_2_cf_exceptionVec_12 ^ toggle_9777_valid_reg;
  assign toggle_9778_clock = clock;
  assign toggle_9778_reset = reset;
  assign toggle_9778_valid = dataBuffer_2_cf_intrVec_1 ^ toggle_9778_valid_reg;
  assign toggle_9779_clock = clock;
  assign toggle_9779_reset = reset;
  assign toggle_9779_valid = dataBuffer_2_cf_intrVec_3 ^ toggle_9779_valid_reg;
  assign toggle_9780_clock = clock;
  assign toggle_9780_reset = reset;
  assign toggle_9780_valid = dataBuffer_2_cf_intrVec_5 ^ toggle_9780_valid_reg;
  assign toggle_9781_clock = clock;
  assign toggle_9781_reset = reset;
  assign toggle_9781_valid = dataBuffer_2_cf_intrVec_7 ^ toggle_9781_valid_reg;
  assign toggle_9782_clock = clock;
  assign toggle_9782_reset = reset;
  assign toggle_9782_valid = dataBuffer_2_cf_intrVec_9 ^ toggle_9782_valid_reg;
  assign toggle_9783_clock = clock;
  assign toggle_9783_reset = reset;
  assign toggle_9783_valid = dataBuffer_2_cf_intrVec_11 ^ toggle_9783_valid_reg;
  assign toggle_9784_clock = clock;
  assign toggle_9784_reset = reset;
  assign toggle_9784_valid = dataBuffer_2_cf_brIdx ^ toggle_9784_valid_reg;
  assign toggle_9788_clock = clock;
  assign toggle_9788_reset = reset;
  assign toggle_9788_valid = dataBuffer_2_cf_crossBoundaryFault ^ toggle_9788_valid_reg;
  assign toggle_9789_clock = clock;
  assign toggle_9789_reset = reset;
  assign toggle_9789_valid = dataBuffer_2_ctrl_src1Type ^ toggle_9789_valid_reg;
  assign toggle_9790_clock = clock;
  assign toggle_9790_reset = reset;
  assign toggle_9790_valid = dataBuffer_2_ctrl_src2Type ^ toggle_9790_valid_reg;
  assign toggle_9791_clock = clock;
  assign toggle_9791_reset = reset;
  assign toggle_9791_valid = dataBuffer_2_ctrl_fuType ^ toggle_9791_valid_reg;
  assign toggle_9794_clock = clock;
  assign toggle_9794_reset = reset;
  assign toggle_9794_valid = dataBuffer_2_ctrl_fuOpType ^ toggle_9794_valid_reg;
  assign toggle_9801_clock = clock;
  assign toggle_9801_reset = reset;
  assign toggle_9801_valid = dataBuffer_2_ctrl_rfSrc1 ^ toggle_9801_valid_reg;
  assign toggle_9806_clock = clock;
  assign toggle_9806_reset = reset;
  assign toggle_9806_valid = dataBuffer_2_ctrl_rfSrc2 ^ toggle_9806_valid_reg;
  assign toggle_9811_clock = clock;
  assign toggle_9811_reset = reset;
  assign toggle_9811_valid = dataBuffer_2_ctrl_rfWen ^ toggle_9811_valid_reg;
  assign toggle_9812_clock = clock;
  assign toggle_9812_reset = reset;
  assign toggle_9812_valid = dataBuffer_2_ctrl_rfDest ^ toggle_9812_valid_reg;
  assign toggle_9817_clock = clock;
  assign toggle_9817_reset = reset;
  assign toggle_9817_valid = dataBuffer_2_ctrl_isNutCoreTrap ^ toggle_9817_valid_reg;
  assign toggle_9818_clock = clock;
  assign toggle_9818_reset = reset;
  assign toggle_9818_valid = dataBuffer_2_data_imm ^ toggle_9818_valid_reg;
  assign toggle_9882_clock = clock;
  assign toggle_9882_reset = reset;
  assign toggle_9882_valid = dataBuffer_3_cf_instr ^ toggle_9882_valid_reg;
  assign toggle_9946_clock = clock;
  assign toggle_9946_reset = reset;
  assign toggle_9946_valid = dataBuffer_3_cf_pc ^ toggle_9946_valid_reg;
  assign toggle_9985_clock = clock;
  assign toggle_9985_reset = reset;
  assign toggle_9985_valid = dataBuffer_3_cf_pnpc ^ toggle_9985_valid_reg;
  assign toggle_10024_clock = clock;
  assign toggle_10024_reset = reset;
  assign toggle_10024_valid = dataBuffer_3_cf_exceptionVec_1 ^ toggle_10024_valid_reg;
  assign toggle_10025_clock = clock;
  assign toggle_10025_reset = reset;
  assign toggle_10025_valid = dataBuffer_3_cf_exceptionVec_2 ^ toggle_10025_valid_reg;
  assign toggle_10026_clock = clock;
  assign toggle_10026_reset = reset;
  assign toggle_10026_valid = dataBuffer_3_cf_exceptionVec_12 ^ toggle_10026_valid_reg;
  assign toggle_10027_clock = clock;
  assign toggle_10027_reset = reset;
  assign toggle_10027_valid = dataBuffer_3_cf_intrVec_1 ^ toggle_10027_valid_reg;
  assign toggle_10028_clock = clock;
  assign toggle_10028_reset = reset;
  assign toggle_10028_valid = dataBuffer_3_cf_intrVec_3 ^ toggle_10028_valid_reg;
  assign toggle_10029_clock = clock;
  assign toggle_10029_reset = reset;
  assign toggle_10029_valid = dataBuffer_3_cf_intrVec_5 ^ toggle_10029_valid_reg;
  assign toggle_10030_clock = clock;
  assign toggle_10030_reset = reset;
  assign toggle_10030_valid = dataBuffer_3_cf_intrVec_7 ^ toggle_10030_valid_reg;
  assign toggle_10031_clock = clock;
  assign toggle_10031_reset = reset;
  assign toggle_10031_valid = dataBuffer_3_cf_intrVec_9 ^ toggle_10031_valid_reg;
  assign toggle_10032_clock = clock;
  assign toggle_10032_reset = reset;
  assign toggle_10032_valid = dataBuffer_3_cf_intrVec_11 ^ toggle_10032_valid_reg;
  assign toggle_10033_clock = clock;
  assign toggle_10033_reset = reset;
  assign toggle_10033_valid = dataBuffer_3_cf_brIdx ^ toggle_10033_valid_reg;
  assign toggle_10037_clock = clock;
  assign toggle_10037_reset = reset;
  assign toggle_10037_valid = dataBuffer_3_cf_crossBoundaryFault ^ toggle_10037_valid_reg;
  assign toggle_10038_clock = clock;
  assign toggle_10038_reset = reset;
  assign toggle_10038_valid = dataBuffer_3_ctrl_src1Type ^ toggle_10038_valid_reg;
  assign toggle_10039_clock = clock;
  assign toggle_10039_reset = reset;
  assign toggle_10039_valid = dataBuffer_3_ctrl_src2Type ^ toggle_10039_valid_reg;
  assign toggle_10040_clock = clock;
  assign toggle_10040_reset = reset;
  assign toggle_10040_valid = dataBuffer_3_ctrl_fuType ^ toggle_10040_valid_reg;
  assign toggle_10043_clock = clock;
  assign toggle_10043_reset = reset;
  assign toggle_10043_valid = dataBuffer_3_ctrl_fuOpType ^ toggle_10043_valid_reg;
  assign toggle_10050_clock = clock;
  assign toggle_10050_reset = reset;
  assign toggle_10050_valid = dataBuffer_3_ctrl_rfSrc1 ^ toggle_10050_valid_reg;
  assign toggle_10055_clock = clock;
  assign toggle_10055_reset = reset;
  assign toggle_10055_valid = dataBuffer_3_ctrl_rfSrc2 ^ toggle_10055_valid_reg;
  assign toggle_10060_clock = clock;
  assign toggle_10060_reset = reset;
  assign toggle_10060_valid = dataBuffer_3_ctrl_rfWen ^ toggle_10060_valid_reg;
  assign toggle_10061_clock = clock;
  assign toggle_10061_reset = reset;
  assign toggle_10061_valid = dataBuffer_3_ctrl_rfDest ^ toggle_10061_valid_reg;
  assign toggle_10066_clock = clock;
  assign toggle_10066_reset = reset;
  assign toggle_10066_valid = dataBuffer_3_ctrl_isNutCoreTrap ^ toggle_10066_valid_reg;
  assign toggle_10067_clock = clock;
  assign toggle_10067_reset = reset;
  assign toggle_10067_valid = dataBuffer_3_data_imm ^ toggle_10067_valid_reg;
  assign toggle_10131_clock = clock;
  assign toggle_10131_reset = reset;
  assign toggle_10131_valid = ringBufferHead ^ toggle_10131_valid_reg;
  assign toggle_10133_clock = clock;
  assign toggle_10133_reset = reset;
  assign toggle_10133_valid = ringBufferTail ^ toggle_10133_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_instr <= _GEN_224;
        end
      end else begin
        dataBuffer_0_cf_instr <= _GEN_224;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_pc <= _GEN_228;
        end
      end else begin
        dataBuffer_0_cf_pc <= _GEN_228;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_pnpc <= _GEN_232;
        end
      end else begin
        dataBuffer_0_cf_pnpc <= _GEN_232;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_exceptionVec_1 <= _GEN_252;
        end
      end else begin
        dataBuffer_0_cf_exceptionVec_1 <= _GEN_252;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_exceptionVec_2 <= _GEN_256;
        end
      end else begin
        dataBuffer_0_cf_exceptionVec_2 <= _GEN_256;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_exceptionVec_12 <= _GEN_296;
        end
      end else begin
        dataBuffer_0_cf_exceptionVec_12 <= _GEN_296;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_1 <= _GEN_316;
        end
      end else begin
        dataBuffer_0_cf_intrVec_1 <= _GEN_316;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_3 <= _GEN_324;
        end
      end else begin
        dataBuffer_0_cf_intrVec_3 <= _GEN_324;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_5 <= _GEN_332;
        end
      end else begin
        dataBuffer_0_cf_intrVec_5 <= _GEN_332;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_7 <= _GEN_340;
        end
      end else begin
        dataBuffer_0_cf_intrVec_7 <= _GEN_340;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_9 <= _GEN_348;
        end
      end else begin
        dataBuffer_0_cf_intrVec_9 <= _GEN_348;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_intrVec_11 <= _GEN_356;
        end
      end else begin
        dataBuffer_0_cf_intrVec_11 <= _GEN_356;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_brIdx <= _GEN_360;
        end
      end else begin
        dataBuffer_0_cf_brIdx <= _GEN_360;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_cf_crossBoundaryFault <= _GEN_368;
        end
      end else begin
        dataBuffer_0_cf_crossBoundaryFault <= _GEN_368;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_src1Type <= _GEN_384;
        end
      end else begin
        dataBuffer_0_ctrl_src1Type <= _GEN_384;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_src2Type <= _GEN_388;
        end
      end else begin
        dataBuffer_0_ctrl_src2Type <= _GEN_388;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_fuType <= _GEN_392;
        end
      end else begin
        dataBuffer_0_ctrl_fuType <= _GEN_392;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_fuOpType <= _GEN_396;
        end
      end else begin
        dataBuffer_0_ctrl_fuOpType <= _GEN_396;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_rfSrc1 <= _GEN_400;
        end
      end else begin
        dataBuffer_0_ctrl_rfSrc1 <= _GEN_400;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_rfSrc2 <= _GEN_404;
        end
      end else begin
        dataBuffer_0_ctrl_rfSrc2 <= _GEN_404;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_rfWen <= _GEN_408;
        end
      end else begin
        dataBuffer_0_ctrl_rfWen <= _GEN_408;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_rfDest <= _GEN_412;
        end
      end else begin
        dataBuffer_0_ctrl_rfDest <= _GEN_412;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_ctrl_isNutCoreTrap <= _GEN_416;
        end
      end else begin
        dataBuffer_0_ctrl_isNutCoreTrap <= _GEN_416;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_0_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h0 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_0_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_0_data_imm <= _GEN_444;
        end
      end else begin
        dataBuffer_0_data_imm <= _GEN_444;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_instr <= _GEN_225;
        end
      end else begin
        dataBuffer_1_cf_instr <= _GEN_225;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_pc <= _GEN_229;
        end
      end else begin
        dataBuffer_1_cf_pc <= _GEN_229;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_pnpc <= _GEN_233;
        end
      end else begin
        dataBuffer_1_cf_pnpc <= _GEN_233;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_exceptionVec_1 <= _GEN_253;
        end
      end else begin
        dataBuffer_1_cf_exceptionVec_1 <= _GEN_253;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_exceptionVec_2 <= _GEN_257;
        end
      end else begin
        dataBuffer_1_cf_exceptionVec_2 <= _GEN_257;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_exceptionVec_12 <= _GEN_297;
        end
      end else begin
        dataBuffer_1_cf_exceptionVec_12 <= _GEN_297;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_1 <= _GEN_317;
        end
      end else begin
        dataBuffer_1_cf_intrVec_1 <= _GEN_317;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_3 <= _GEN_325;
        end
      end else begin
        dataBuffer_1_cf_intrVec_3 <= _GEN_325;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_5 <= _GEN_333;
        end
      end else begin
        dataBuffer_1_cf_intrVec_5 <= _GEN_333;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_7 <= _GEN_341;
        end
      end else begin
        dataBuffer_1_cf_intrVec_7 <= _GEN_341;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_9 <= _GEN_349;
        end
      end else begin
        dataBuffer_1_cf_intrVec_9 <= _GEN_349;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_intrVec_11 <= _GEN_357;
        end
      end else begin
        dataBuffer_1_cf_intrVec_11 <= _GEN_357;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_brIdx <= _GEN_361;
        end
      end else begin
        dataBuffer_1_cf_brIdx <= _GEN_361;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_cf_crossBoundaryFault <= _GEN_369;
        end
      end else begin
        dataBuffer_1_cf_crossBoundaryFault <= _GEN_369;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_src1Type <= _GEN_385;
        end
      end else begin
        dataBuffer_1_ctrl_src1Type <= _GEN_385;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_src2Type <= _GEN_389;
        end
      end else begin
        dataBuffer_1_ctrl_src2Type <= _GEN_389;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_fuType <= _GEN_393;
        end
      end else begin
        dataBuffer_1_ctrl_fuType <= _GEN_393;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_fuOpType <= _GEN_397;
        end
      end else begin
        dataBuffer_1_ctrl_fuOpType <= _GEN_397;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_rfSrc1 <= _GEN_401;
        end
      end else begin
        dataBuffer_1_ctrl_rfSrc1 <= _GEN_401;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_rfSrc2 <= _GEN_405;
        end
      end else begin
        dataBuffer_1_ctrl_rfSrc2 <= _GEN_405;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_rfWen <= _GEN_409;
        end
      end else begin
        dataBuffer_1_ctrl_rfWen <= _GEN_409;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_rfDest <= _GEN_413;
        end
      end else begin
        dataBuffer_1_ctrl_rfDest <= _GEN_413;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_ctrl_isNutCoreTrap <= _GEN_417;
        end
      end else begin
        dataBuffer_1_ctrl_isNutCoreTrap <= _GEN_417;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_1_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h1 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_1_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_1_data_imm <= _GEN_445;
        end
      end else begin
        dataBuffer_1_data_imm <= _GEN_445;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_instr <= _GEN_226;
        end
      end else begin
        dataBuffer_2_cf_instr <= _GEN_226;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_pc <= _GEN_230;
        end
      end else begin
        dataBuffer_2_cf_pc <= _GEN_230;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_pnpc <= _GEN_234;
        end
      end else begin
        dataBuffer_2_cf_pnpc <= _GEN_234;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_exceptionVec_1 <= _GEN_254;
        end
      end else begin
        dataBuffer_2_cf_exceptionVec_1 <= _GEN_254;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_exceptionVec_2 <= _GEN_258;
        end
      end else begin
        dataBuffer_2_cf_exceptionVec_2 <= _GEN_258;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_exceptionVec_12 <= _GEN_298;
        end
      end else begin
        dataBuffer_2_cf_exceptionVec_12 <= _GEN_298;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_1 <= _GEN_318;
        end
      end else begin
        dataBuffer_2_cf_intrVec_1 <= _GEN_318;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_3 <= _GEN_326;
        end
      end else begin
        dataBuffer_2_cf_intrVec_3 <= _GEN_326;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_5 <= _GEN_334;
        end
      end else begin
        dataBuffer_2_cf_intrVec_5 <= _GEN_334;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_7 <= _GEN_342;
        end
      end else begin
        dataBuffer_2_cf_intrVec_7 <= _GEN_342;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_9 <= _GEN_350;
        end
      end else begin
        dataBuffer_2_cf_intrVec_9 <= _GEN_350;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_intrVec_11 <= _GEN_358;
        end
      end else begin
        dataBuffer_2_cf_intrVec_11 <= _GEN_358;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_brIdx <= _GEN_362;
        end
      end else begin
        dataBuffer_2_cf_brIdx <= _GEN_362;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_cf_crossBoundaryFault <= _GEN_370;
        end
      end else begin
        dataBuffer_2_cf_crossBoundaryFault <= _GEN_370;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_src1Type <= _GEN_386;
        end
      end else begin
        dataBuffer_2_ctrl_src1Type <= _GEN_386;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_src2Type <= _GEN_390;
        end
      end else begin
        dataBuffer_2_ctrl_src2Type <= _GEN_390;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_fuType <= _GEN_394;
        end
      end else begin
        dataBuffer_2_ctrl_fuType <= _GEN_394;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_fuOpType <= _GEN_398;
        end
      end else begin
        dataBuffer_2_ctrl_fuOpType <= _GEN_398;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_rfSrc1 <= _GEN_402;
        end
      end else begin
        dataBuffer_2_ctrl_rfSrc1 <= _GEN_402;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_rfSrc2 <= _GEN_406;
        end
      end else begin
        dataBuffer_2_ctrl_rfSrc2 <= _GEN_406;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_rfWen <= _GEN_410;
        end
      end else begin
        dataBuffer_2_ctrl_rfWen <= _GEN_410;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_rfDest <= _GEN_414;
        end
      end else begin
        dataBuffer_2_ctrl_rfDest <= _GEN_414;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_ctrl_isNutCoreTrap <= _GEN_418;
        end
      end else begin
        dataBuffer_2_ctrl_isNutCoreTrap <= _GEN_418;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_2_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h2 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_2_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_2_data_imm <= _GEN_446;
        end
      end else begin
        dataBuffer_2_data_imm <= _GEN_446;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_instr <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_instr <= _GEN_227;
        end
      end else begin
        dataBuffer_3_cf_instr <= _GEN_227;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_pc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_pc <= _GEN_231;
        end
      end else begin
        dataBuffer_3_cf_pc <= _GEN_231;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_pnpc <= 39'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_pnpc <= _GEN_235;
        end
      end else begin
        dataBuffer_3_cf_pnpc <= _GEN_235;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_exceptionVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_exceptionVec_1 <= _GEN_255;
        end
      end else begin
        dataBuffer_3_cf_exceptionVec_1 <= _GEN_255;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_exceptionVec_2 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_exceptionVec_2 <= _GEN_259;
        end
      end else begin
        dataBuffer_3_cf_exceptionVec_2 <= _GEN_259;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_exceptionVec_12 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_exceptionVec_12 <= _GEN_299;
        end
      end else begin
        dataBuffer_3_cf_exceptionVec_12 <= _GEN_299;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_1 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_1 <= _GEN_319;
        end
      end else begin
        dataBuffer_3_cf_intrVec_1 <= _GEN_319;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_3 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_3 <= _GEN_327;
        end
      end else begin
        dataBuffer_3_cf_intrVec_3 <= _GEN_327;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_5 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_5 <= _GEN_335;
        end
      end else begin
        dataBuffer_3_cf_intrVec_5 <= _GEN_335;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_7 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_7 <= _GEN_343;
        end
      end else begin
        dataBuffer_3_cf_intrVec_7 <= _GEN_343;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_9 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_9 <= _GEN_351;
        end
      end else begin
        dataBuffer_3_cf_intrVec_9 <= _GEN_351;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_intrVec_11 <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_intrVec_11 <= _GEN_359;
        end
      end else begin
        dataBuffer_3_cf_intrVec_11 <= _GEN_359;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_brIdx <= 4'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_brIdx <= _GEN_363;
        end
      end else begin
        dataBuffer_3_cf_brIdx <= _GEN_363;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_cf_crossBoundaryFault <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_cf_crossBoundaryFault <= _GEN_371;
        end
      end else begin
        dataBuffer_3_cf_crossBoundaryFault <= _GEN_371;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_src1Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_src1Type <= _GEN_387;
        end
      end else begin
        dataBuffer_3_ctrl_src1Type <= _GEN_387;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_src2Type <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_src2Type <= _GEN_391;
        end
      end else begin
        dataBuffer_3_ctrl_src2Type <= _GEN_391;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_fuType <= 3'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_fuType <= _GEN_395;
        end
      end else begin
        dataBuffer_3_ctrl_fuType <= _GEN_395;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_fuOpType <= 7'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_fuOpType <= _GEN_399;
        end
      end else begin
        dataBuffer_3_ctrl_fuOpType <= _GEN_399;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_rfSrc1 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_rfSrc1 <= _GEN_403;
        end
      end else begin
        dataBuffer_3_ctrl_rfSrc1 <= _GEN_403;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_rfSrc2 <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_rfSrc2 <= _GEN_407;
        end
      end else begin
        dataBuffer_3_ctrl_rfSrc2 <= _GEN_407;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_rfWen <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_rfWen <= _GEN_411;
        end
      end else begin
        dataBuffer_3_ctrl_rfWen <= _GEN_411;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_rfDest <= 5'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_rfDest <= _GEN_415;
        end
      end else begin
        dataBuffer_3_ctrl_rfDest <= _GEN_415;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_ctrl_isNutCoreTrap <= 1'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_ctrl_isNutCoreTrap <= _GEN_419;
        end
      end else begin
        dataBuffer_3_ctrl_isNutCoreTrap <= _GEN_419;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 29:29]
      dataBuffer_3_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      if (enqueueFire_1) begin // @[src/main/scala/utils/PipelineVector.scala 46:29]
        if (2'h3 == _T_4) begin // @[src/main/scala/utils/PipelineVector.scala 46:63]
          dataBuffer_3_data_imm <= 64'h0; // @[src/main/scala/utils/PipelineVector.scala 46:63]
        end else begin
          dataBuffer_3_data_imm <= _GEN_447;
        end
      end else begin
        dataBuffer_3_data_imm <= _GEN_447;
      end
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 30:33]
      ringBufferHead <= 2'h0; // @[src/main/scala/utils/PipelineVector.scala 30:33]
    end else if (frontend_io_flushVec[1]) begin // @[src/main/scala/utils/PipelineVector.scala 71:16]
      ringBufferHead <= 2'h0; // @[src/main/scala/utils/PipelineVector.scala 72:24]
    end else if (wen) begin // @[src/main/scala/utils/PipelineVector.scala 44:14]
      ringBufferHead <= _ringBufferHead_T_1; // @[src/main/scala/utils/PipelineVector.scala 47:24]
    end
    if (reset) begin // @[src/main/scala/utils/PipelineVector.scala 31:33]
      ringBufferTail <= 2'h0; // @[src/main/scala/utils/PipelineVector.scala 31:33]
    end else if (frontend_io_flushVec[1]) begin // @[src/main/scala/utils/PipelineVector.scala 71:16]
      ringBufferTail <= 2'h0; // @[src/main/scala/utils/PipelineVector.scala 73:24]
    end else if (dequeueFire) begin // @[src/main/scala/utils/PipelineVector.scala 66:22]
      ringBufferTail <= _ringBufferTail_T_1; // @[src/main/scala/utils/PipelineVector.scala 67:24]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    dataBuffer_0_cf_instr_p <= dataBuffer_0_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9135_valid_reg <= dataBuffer_0_cf_instr;
    dataBuffer_0_cf_pc_p <= dataBuffer_0_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9199_valid_reg <= dataBuffer_0_cf_pc;
    dataBuffer_0_cf_pnpc_p <= dataBuffer_0_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9238_valid_reg <= dataBuffer_0_cf_pnpc;
    dataBuffer_0_cf_exceptionVec_1_p <= dataBuffer_0_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9277_valid_reg <= dataBuffer_0_cf_exceptionVec_1;
    dataBuffer_0_cf_exceptionVec_2_p <= dataBuffer_0_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9278_valid_reg <= dataBuffer_0_cf_exceptionVec_2;
    dataBuffer_0_cf_exceptionVec_12_p <= dataBuffer_0_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9279_valid_reg <= dataBuffer_0_cf_exceptionVec_12;
    dataBuffer_0_cf_intrVec_1_p <= dataBuffer_0_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9280_valid_reg <= dataBuffer_0_cf_intrVec_1;
    dataBuffer_0_cf_intrVec_3_p <= dataBuffer_0_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9281_valid_reg <= dataBuffer_0_cf_intrVec_3;
    dataBuffer_0_cf_intrVec_5_p <= dataBuffer_0_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9282_valid_reg <= dataBuffer_0_cf_intrVec_5;
    dataBuffer_0_cf_intrVec_7_p <= dataBuffer_0_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9283_valid_reg <= dataBuffer_0_cf_intrVec_7;
    dataBuffer_0_cf_intrVec_9_p <= dataBuffer_0_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9284_valid_reg <= dataBuffer_0_cf_intrVec_9;
    dataBuffer_0_cf_intrVec_11_p <= dataBuffer_0_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9285_valid_reg <= dataBuffer_0_cf_intrVec_11;
    dataBuffer_0_cf_brIdx_p <= dataBuffer_0_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9286_valid_reg <= dataBuffer_0_cf_brIdx;
    dataBuffer_0_cf_crossBoundaryFault_p <= dataBuffer_0_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9290_valid_reg <= dataBuffer_0_cf_crossBoundaryFault;
    dataBuffer_0_ctrl_src1Type_p <= dataBuffer_0_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9291_valid_reg <= dataBuffer_0_ctrl_src1Type;
    dataBuffer_0_ctrl_src2Type_p <= dataBuffer_0_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9292_valid_reg <= dataBuffer_0_ctrl_src2Type;
    dataBuffer_0_ctrl_fuType_p <= dataBuffer_0_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9293_valid_reg <= dataBuffer_0_ctrl_fuType;
    dataBuffer_0_ctrl_fuOpType_p <= dataBuffer_0_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9296_valid_reg <= dataBuffer_0_ctrl_fuOpType;
    dataBuffer_0_ctrl_rfSrc1_p <= dataBuffer_0_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9303_valid_reg <= dataBuffer_0_ctrl_rfSrc1;
    dataBuffer_0_ctrl_rfSrc2_p <= dataBuffer_0_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9308_valid_reg <= dataBuffer_0_ctrl_rfSrc2;
    dataBuffer_0_ctrl_rfWen_p <= dataBuffer_0_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9313_valid_reg <= dataBuffer_0_ctrl_rfWen;
    dataBuffer_0_ctrl_rfDest_p <= dataBuffer_0_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9314_valid_reg <= dataBuffer_0_ctrl_rfDest;
    dataBuffer_0_ctrl_isNutCoreTrap_p <= dataBuffer_0_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9319_valid_reg <= dataBuffer_0_ctrl_isNutCoreTrap;
    dataBuffer_0_data_imm_p <= dataBuffer_0_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9320_valid_reg <= dataBuffer_0_data_imm;
    dataBuffer_1_cf_instr_p <= dataBuffer_1_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9384_valid_reg <= dataBuffer_1_cf_instr;
    dataBuffer_1_cf_pc_p <= dataBuffer_1_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9448_valid_reg <= dataBuffer_1_cf_pc;
    dataBuffer_1_cf_pnpc_p <= dataBuffer_1_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9487_valid_reg <= dataBuffer_1_cf_pnpc;
    dataBuffer_1_cf_exceptionVec_1_p <= dataBuffer_1_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9526_valid_reg <= dataBuffer_1_cf_exceptionVec_1;
    dataBuffer_1_cf_exceptionVec_2_p <= dataBuffer_1_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9527_valid_reg <= dataBuffer_1_cf_exceptionVec_2;
    dataBuffer_1_cf_exceptionVec_12_p <= dataBuffer_1_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9528_valid_reg <= dataBuffer_1_cf_exceptionVec_12;
    dataBuffer_1_cf_intrVec_1_p <= dataBuffer_1_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9529_valid_reg <= dataBuffer_1_cf_intrVec_1;
    dataBuffer_1_cf_intrVec_3_p <= dataBuffer_1_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9530_valid_reg <= dataBuffer_1_cf_intrVec_3;
    dataBuffer_1_cf_intrVec_5_p <= dataBuffer_1_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9531_valid_reg <= dataBuffer_1_cf_intrVec_5;
    dataBuffer_1_cf_intrVec_7_p <= dataBuffer_1_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9532_valid_reg <= dataBuffer_1_cf_intrVec_7;
    dataBuffer_1_cf_intrVec_9_p <= dataBuffer_1_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9533_valid_reg <= dataBuffer_1_cf_intrVec_9;
    dataBuffer_1_cf_intrVec_11_p <= dataBuffer_1_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9534_valid_reg <= dataBuffer_1_cf_intrVec_11;
    dataBuffer_1_cf_brIdx_p <= dataBuffer_1_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9535_valid_reg <= dataBuffer_1_cf_brIdx;
    dataBuffer_1_cf_crossBoundaryFault_p <= dataBuffer_1_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9539_valid_reg <= dataBuffer_1_cf_crossBoundaryFault;
    dataBuffer_1_ctrl_src1Type_p <= dataBuffer_1_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9540_valid_reg <= dataBuffer_1_ctrl_src1Type;
    dataBuffer_1_ctrl_src2Type_p <= dataBuffer_1_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9541_valid_reg <= dataBuffer_1_ctrl_src2Type;
    dataBuffer_1_ctrl_fuType_p <= dataBuffer_1_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9542_valid_reg <= dataBuffer_1_ctrl_fuType;
    dataBuffer_1_ctrl_fuOpType_p <= dataBuffer_1_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9545_valid_reg <= dataBuffer_1_ctrl_fuOpType;
    dataBuffer_1_ctrl_rfSrc1_p <= dataBuffer_1_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9552_valid_reg <= dataBuffer_1_ctrl_rfSrc1;
    dataBuffer_1_ctrl_rfSrc2_p <= dataBuffer_1_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9557_valid_reg <= dataBuffer_1_ctrl_rfSrc2;
    dataBuffer_1_ctrl_rfWen_p <= dataBuffer_1_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9562_valid_reg <= dataBuffer_1_ctrl_rfWen;
    dataBuffer_1_ctrl_rfDest_p <= dataBuffer_1_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9563_valid_reg <= dataBuffer_1_ctrl_rfDest;
    dataBuffer_1_ctrl_isNutCoreTrap_p <= dataBuffer_1_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9568_valid_reg <= dataBuffer_1_ctrl_isNutCoreTrap;
    dataBuffer_1_data_imm_p <= dataBuffer_1_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9569_valid_reg <= dataBuffer_1_data_imm;
    dataBuffer_2_cf_instr_p <= dataBuffer_2_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9633_valid_reg <= dataBuffer_2_cf_instr;
    dataBuffer_2_cf_pc_p <= dataBuffer_2_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9697_valid_reg <= dataBuffer_2_cf_pc;
    dataBuffer_2_cf_pnpc_p <= dataBuffer_2_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9736_valid_reg <= dataBuffer_2_cf_pnpc;
    dataBuffer_2_cf_exceptionVec_1_p <= dataBuffer_2_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9775_valid_reg <= dataBuffer_2_cf_exceptionVec_1;
    dataBuffer_2_cf_exceptionVec_2_p <= dataBuffer_2_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9776_valid_reg <= dataBuffer_2_cf_exceptionVec_2;
    dataBuffer_2_cf_exceptionVec_12_p <= dataBuffer_2_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9777_valid_reg <= dataBuffer_2_cf_exceptionVec_12;
    dataBuffer_2_cf_intrVec_1_p <= dataBuffer_2_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9778_valid_reg <= dataBuffer_2_cf_intrVec_1;
    dataBuffer_2_cf_intrVec_3_p <= dataBuffer_2_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9779_valid_reg <= dataBuffer_2_cf_intrVec_3;
    dataBuffer_2_cf_intrVec_5_p <= dataBuffer_2_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9780_valid_reg <= dataBuffer_2_cf_intrVec_5;
    dataBuffer_2_cf_intrVec_7_p <= dataBuffer_2_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9781_valid_reg <= dataBuffer_2_cf_intrVec_7;
    dataBuffer_2_cf_intrVec_9_p <= dataBuffer_2_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9782_valid_reg <= dataBuffer_2_cf_intrVec_9;
    dataBuffer_2_cf_intrVec_11_p <= dataBuffer_2_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9783_valid_reg <= dataBuffer_2_cf_intrVec_11;
    dataBuffer_2_cf_brIdx_p <= dataBuffer_2_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9784_valid_reg <= dataBuffer_2_cf_brIdx;
    dataBuffer_2_cf_crossBoundaryFault_p <= dataBuffer_2_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9788_valid_reg <= dataBuffer_2_cf_crossBoundaryFault;
    dataBuffer_2_ctrl_src1Type_p <= dataBuffer_2_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9789_valid_reg <= dataBuffer_2_ctrl_src1Type;
    dataBuffer_2_ctrl_src2Type_p <= dataBuffer_2_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9790_valid_reg <= dataBuffer_2_ctrl_src2Type;
    dataBuffer_2_ctrl_fuType_p <= dataBuffer_2_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9791_valid_reg <= dataBuffer_2_ctrl_fuType;
    dataBuffer_2_ctrl_fuOpType_p <= dataBuffer_2_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9794_valid_reg <= dataBuffer_2_ctrl_fuOpType;
    dataBuffer_2_ctrl_rfSrc1_p <= dataBuffer_2_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9801_valid_reg <= dataBuffer_2_ctrl_rfSrc1;
    dataBuffer_2_ctrl_rfSrc2_p <= dataBuffer_2_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9806_valid_reg <= dataBuffer_2_ctrl_rfSrc2;
    dataBuffer_2_ctrl_rfWen_p <= dataBuffer_2_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9811_valid_reg <= dataBuffer_2_ctrl_rfWen;
    dataBuffer_2_ctrl_rfDest_p <= dataBuffer_2_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9812_valid_reg <= dataBuffer_2_ctrl_rfDest;
    dataBuffer_2_ctrl_isNutCoreTrap_p <= dataBuffer_2_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9817_valid_reg <= dataBuffer_2_ctrl_isNutCoreTrap;
    dataBuffer_2_data_imm_p <= dataBuffer_2_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9818_valid_reg <= dataBuffer_2_data_imm;
    dataBuffer_3_cf_instr_p <= dataBuffer_3_cf_instr; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9882_valid_reg <= dataBuffer_3_cf_instr;
    dataBuffer_3_cf_pc_p <= dataBuffer_3_cf_pc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9946_valid_reg <= dataBuffer_3_cf_pc;
    dataBuffer_3_cf_pnpc_p <= dataBuffer_3_cf_pnpc; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_9985_valid_reg <= dataBuffer_3_cf_pnpc;
    dataBuffer_3_cf_exceptionVec_1_p <= dataBuffer_3_cf_exceptionVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10024_valid_reg <= dataBuffer_3_cf_exceptionVec_1;
    dataBuffer_3_cf_exceptionVec_2_p <= dataBuffer_3_cf_exceptionVec_2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10025_valid_reg <= dataBuffer_3_cf_exceptionVec_2;
    dataBuffer_3_cf_exceptionVec_12_p <= dataBuffer_3_cf_exceptionVec_12; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10026_valid_reg <= dataBuffer_3_cf_exceptionVec_12;
    dataBuffer_3_cf_intrVec_1_p <= dataBuffer_3_cf_intrVec_1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10027_valid_reg <= dataBuffer_3_cf_intrVec_1;
    dataBuffer_3_cf_intrVec_3_p <= dataBuffer_3_cf_intrVec_3; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10028_valid_reg <= dataBuffer_3_cf_intrVec_3;
    dataBuffer_3_cf_intrVec_5_p <= dataBuffer_3_cf_intrVec_5; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10029_valid_reg <= dataBuffer_3_cf_intrVec_5;
    dataBuffer_3_cf_intrVec_7_p <= dataBuffer_3_cf_intrVec_7; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10030_valid_reg <= dataBuffer_3_cf_intrVec_7;
    dataBuffer_3_cf_intrVec_9_p <= dataBuffer_3_cf_intrVec_9; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10031_valid_reg <= dataBuffer_3_cf_intrVec_9;
    dataBuffer_3_cf_intrVec_11_p <= dataBuffer_3_cf_intrVec_11; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10032_valid_reg <= dataBuffer_3_cf_intrVec_11;
    dataBuffer_3_cf_brIdx_p <= dataBuffer_3_cf_brIdx; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10033_valid_reg <= dataBuffer_3_cf_brIdx;
    dataBuffer_3_cf_crossBoundaryFault_p <= dataBuffer_3_cf_crossBoundaryFault; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10037_valid_reg <= dataBuffer_3_cf_crossBoundaryFault;
    dataBuffer_3_ctrl_src1Type_p <= dataBuffer_3_ctrl_src1Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10038_valid_reg <= dataBuffer_3_ctrl_src1Type;
    dataBuffer_3_ctrl_src2Type_p <= dataBuffer_3_ctrl_src2Type; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10039_valid_reg <= dataBuffer_3_ctrl_src2Type;
    dataBuffer_3_ctrl_fuType_p <= dataBuffer_3_ctrl_fuType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10040_valid_reg <= dataBuffer_3_ctrl_fuType;
    dataBuffer_3_ctrl_fuOpType_p <= dataBuffer_3_ctrl_fuOpType; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10043_valid_reg <= dataBuffer_3_ctrl_fuOpType;
    dataBuffer_3_ctrl_rfSrc1_p <= dataBuffer_3_ctrl_rfSrc1; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10050_valid_reg <= dataBuffer_3_ctrl_rfSrc1;
    dataBuffer_3_ctrl_rfSrc2_p <= dataBuffer_3_ctrl_rfSrc2; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10055_valid_reg <= dataBuffer_3_ctrl_rfSrc2;
    dataBuffer_3_ctrl_rfWen_p <= dataBuffer_3_ctrl_rfWen; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10060_valid_reg <= dataBuffer_3_ctrl_rfWen;
    dataBuffer_3_ctrl_rfDest_p <= dataBuffer_3_ctrl_rfDest; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10061_valid_reg <= dataBuffer_3_ctrl_rfDest;
    dataBuffer_3_ctrl_isNutCoreTrap_p <= dataBuffer_3_ctrl_isNutCoreTrap; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10066_valid_reg <= dataBuffer_3_ctrl_isNutCoreTrap;
    dataBuffer_3_data_imm_p <= dataBuffer_3_data_imm; // @[src/main/scala/utils/PipelineVector.scala 29:29]
    toggle_10067_valid_reg <= dataBuffer_3_data_imm;
    ringBufferHead_p <= ringBufferHead; // @[src/main/scala/utils/PipelineVector.scala 30:33]
    toggle_10131_valid_reg <= ringBufferHead;
    ringBufferTail_p <= ringBufferTail; // @[src/main/scala/utils/PipelineVector.scala 31:33]
    toggle_10133_valid_reg <= ringBufferTail;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  dataBuffer_0_cf_instr = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  dataBuffer_0_cf_pc = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  dataBuffer_0_cf_pnpc = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  dataBuffer_0_cf_exceptionVec_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  dataBuffer_0_cf_exceptionVec_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  dataBuffer_0_cf_exceptionVec_12 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_5 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_7 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_9 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  dataBuffer_0_cf_brIdx = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  dataBuffer_0_cf_crossBoundaryFault = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  dataBuffer_0_ctrl_src1Type = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  dataBuffer_0_ctrl_src2Type = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  dataBuffer_0_ctrl_fuType = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  dataBuffer_0_ctrl_fuOpType = _RAND_17[6:0];
  _RAND_18 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfSrc1 = _RAND_18[4:0];
  _RAND_19 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfSrc2 = _RAND_19[4:0];
  _RAND_20 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfWen = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfDest = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  dataBuffer_0_ctrl_isNutCoreTrap = _RAND_22[0:0];
  _RAND_23 = {2{`RANDOM}};
  dataBuffer_0_data_imm = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  dataBuffer_1_cf_instr = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  dataBuffer_1_cf_pc = _RAND_25[38:0];
  _RAND_26 = {2{`RANDOM}};
  dataBuffer_1_cf_pnpc = _RAND_26[38:0];
  _RAND_27 = {1{`RANDOM}};
  dataBuffer_1_cf_exceptionVec_1 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  dataBuffer_1_cf_exceptionVec_2 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  dataBuffer_1_cf_exceptionVec_12 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_1 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_3 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_5 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_7 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_9 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_11 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  dataBuffer_1_cf_brIdx = _RAND_36[3:0];
  _RAND_37 = {1{`RANDOM}};
  dataBuffer_1_cf_crossBoundaryFault = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  dataBuffer_1_ctrl_src1Type = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  dataBuffer_1_ctrl_src2Type = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  dataBuffer_1_ctrl_fuType = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  dataBuffer_1_ctrl_fuOpType = _RAND_41[6:0];
  _RAND_42 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfSrc1 = _RAND_42[4:0];
  _RAND_43 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfSrc2 = _RAND_43[4:0];
  _RAND_44 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfWen = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfDest = _RAND_45[4:0];
  _RAND_46 = {1{`RANDOM}};
  dataBuffer_1_ctrl_isNutCoreTrap = _RAND_46[0:0];
  _RAND_47 = {2{`RANDOM}};
  dataBuffer_1_data_imm = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  dataBuffer_2_cf_instr = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  dataBuffer_2_cf_pc = _RAND_49[38:0];
  _RAND_50 = {2{`RANDOM}};
  dataBuffer_2_cf_pnpc = _RAND_50[38:0];
  _RAND_51 = {1{`RANDOM}};
  dataBuffer_2_cf_exceptionVec_1 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  dataBuffer_2_cf_exceptionVec_2 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  dataBuffer_2_cf_exceptionVec_12 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_1 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_3 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_5 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_7 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_9 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_11 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  dataBuffer_2_cf_brIdx = _RAND_60[3:0];
  _RAND_61 = {1{`RANDOM}};
  dataBuffer_2_cf_crossBoundaryFault = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  dataBuffer_2_ctrl_src1Type = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  dataBuffer_2_ctrl_src2Type = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  dataBuffer_2_ctrl_fuType = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  dataBuffer_2_ctrl_fuOpType = _RAND_65[6:0];
  _RAND_66 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfSrc1 = _RAND_66[4:0];
  _RAND_67 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfSrc2 = _RAND_67[4:0];
  _RAND_68 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfWen = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfDest = _RAND_69[4:0];
  _RAND_70 = {1{`RANDOM}};
  dataBuffer_2_ctrl_isNutCoreTrap = _RAND_70[0:0];
  _RAND_71 = {2{`RANDOM}};
  dataBuffer_2_data_imm = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  dataBuffer_3_cf_instr = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  dataBuffer_3_cf_pc = _RAND_73[38:0];
  _RAND_74 = {2{`RANDOM}};
  dataBuffer_3_cf_pnpc = _RAND_74[38:0];
  _RAND_75 = {1{`RANDOM}};
  dataBuffer_3_cf_exceptionVec_1 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  dataBuffer_3_cf_exceptionVec_2 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  dataBuffer_3_cf_exceptionVec_12 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_1 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_3 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_5 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_7 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_9 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_11 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  dataBuffer_3_cf_brIdx = _RAND_84[3:0];
  _RAND_85 = {1{`RANDOM}};
  dataBuffer_3_cf_crossBoundaryFault = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  dataBuffer_3_ctrl_src1Type = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  dataBuffer_3_ctrl_src2Type = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  dataBuffer_3_ctrl_fuType = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  dataBuffer_3_ctrl_fuOpType = _RAND_89[6:0];
  _RAND_90 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfSrc1 = _RAND_90[4:0];
  _RAND_91 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfSrc2 = _RAND_91[4:0];
  _RAND_92 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfWen = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfDest = _RAND_93[4:0];
  _RAND_94 = {1{`RANDOM}};
  dataBuffer_3_ctrl_isNutCoreTrap = _RAND_94[0:0];
  _RAND_95 = {2{`RANDOM}};
  dataBuffer_3_data_imm = _RAND_95[63:0];
  _RAND_96 = {1{`RANDOM}};
  ringBufferHead = _RAND_96[1:0];
  _RAND_97 = {1{`RANDOM}};
  ringBufferTail = _RAND_97[1:0];
  _RAND_98 = {2{`RANDOM}};
  dataBuffer_0_cf_instr_p = _RAND_98[63:0];
  _RAND_99 = {2{`RANDOM}};
  toggle_9135_valid_reg = _RAND_99[63:0];
  _RAND_100 = {2{`RANDOM}};
  dataBuffer_0_cf_pc_p = _RAND_100[38:0];
  _RAND_101 = {2{`RANDOM}};
  toggle_9199_valid_reg = _RAND_101[38:0];
  _RAND_102 = {2{`RANDOM}};
  dataBuffer_0_cf_pnpc_p = _RAND_102[38:0];
  _RAND_103 = {2{`RANDOM}};
  toggle_9238_valid_reg = _RAND_103[38:0];
  _RAND_104 = {1{`RANDOM}};
  dataBuffer_0_cf_exceptionVec_1_p = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  toggle_9277_valid_reg = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  dataBuffer_0_cf_exceptionVec_2_p = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  toggle_9278_valid_reg = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  dataBuffer_0_cf_exceptionVec_12_p = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  toggle_9279_valid_reg = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_1_p = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  toggle_9280_valid_reg = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_3_p = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  toggle_9281_valid_reg = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_5_p = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  toggle_9282_valid_reg = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_7_p = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  toggle_9283_valid_reg = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_9_p = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  toggle_9284_valid_reg = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  dataBuffer_0_cf_intrVec_11_p = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  toggle_9285_valid_reg = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  dataBuffer_0_cf_brIdx_p = _RAND_122[3:0];
  _RAND_123 = {1{`RANDOM}};
  toggle_9286_valid_reg = _RAND_123[3:0];
  _RAND_124 = {1{`RANDOM}};
  dataBuffer_0_cf_crossBoundaryFault_p = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  toggle_9290_valid_reg = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  dataBuffer_0_ctrl_src1Type_p = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  toggle_9291_valid_reg = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  dataBuffer_0_ctrl_src2Type_p = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  toggle_9292_valid_reg = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  dataBuffer_0_ctrl_fuType_p = _RAND_130[2:0];
  _RAND_131 = {1{`RANDOM}};
  toggle_9293_valid_reg = _RAND_131[2:0];
  _RAND_132 = {1{`RANDOM}};
  dataBuffer_0_ctrl_fuOpType_p = _RAND_132[6:0];
  _RAND_133 = {1{`RANDOM}};
  toggle_9296_valid_reg = _RAND_133[6:0];
  _RAND_134 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfSrc1_p = _RAND_134[4:0];
  _RAND_135 = {1{`RANDOM}};
  toggle_9303_valid_reg = _RAND_135[4:0];
  _RAND_136 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfSrc2_p = _RAND_136[4:0];
  _RAND_137 = {1{`RANDOM}};
  toggle_9308_valid_reg = _RAND_137[4:0];
  _RAND_138 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfWen_p = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  toggle_9313_valid_reg = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  dataBuffer_0_ctrl_rfDest_p = _RAND_140[4:0];
  _RAND_141 = {1{`RANDOM}};
  toggle_9314_valid_reg = _RAND_141[4:0];
  _RAND_142 = {1{`RANDOM}};
  dataBuffer_0_ctrl_isNutCoreTrap_p = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  toggle_9319_valid_reg = _RAND_143[0:0];
  _RAND_144 = {2{`RANDOM}};
  dataBuffer_0_data_imm_p = _RAND_144[63:0];
  _RAND_145 = {2{`RANDOM}};
  toggle_9320_valid_reg = _RAND_145[63:0];
  _RAND_146 = {2{`RANDOM}};
  dataBuffer_1_cf_instr_p = _RAND_146[63:0];
  _RAND_147 = {2{`RANDOM}};
  toggle_9384_valid_reg = _RAND_147[63:0];
  _RAND_148 = {2{`RANDOM}};
  dataBuffer_1_cf_pc_p = _RAND_148[38:0];
  _RAND_149 = {2{`RANDOM}};
  toggle_9448_valid_reg = _RAND_149[38:0];
  _RAND_150 = {2{`RANDOM}};
  dataBuffer_1_cf_pnpc_p = _RAND_150[38:0];
  _RAND_151 = {2{`RANDOM}};
  toggle_9487_valid_reg = _RAND_151[38:0];
  _RAND_152 = {1{`RANDOM}};
  dataBuffer_1_cf_exceptionVec_1_p = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  toggle_9526_valid_reg = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  dataBuffer_1_cf_exceptionVec_2_p = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  toggle_9527_valid_reg = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  dataBuffer_1_cf_exceptionVec_12_p = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  toggle_9528_valid_reg = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_1_p = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  toggle_9529_valid_reg = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_3_p = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  toggle_9530_valid_reg = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_5_p = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  toggle_9531_valid_reg = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_7_p = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  toggle_9532_valid_reg = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_9_p = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  toggle_9533_valid_reg = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  dataBuffer_1_cf_intrVec_11_p = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  toggle_9534_valid_reg = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  dataBuffer_1_cf_brIdx_p = _RAND_170[3:0];
  _RAND_171 = {1{`RANDOM}};
  toggle_9535_valid_reg = _RAND_171[3:0];
  _RAND_172 = {1{`RANDOM}};
  dataBuffer_1_cf_crossBoundaryFault_p = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  toggle_9539_valid_reg = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  dataBuffer_1_ctrl_src1Type_p = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  toggle_9540_valid_reg = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  dataBuffer_1_ctrl_src2Type_p = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  toggle_9541_valid_reg = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  dataBuffer_1_ctrl_fuType_p = _RAND_178[2:0];
  _RAND_179 = {1{`RANDOM}};
  toggle_9542_valid_reg = _RAND_179[2:0];
  _RAND_180 = {1{`RANDOM}};
  dataBuffer_1_ctrl_fuOpType_p = _RAND_180[6:0];
  _RAND_181 = {1{`RANDOM}};
  toggle_9545_valid_reg = _RAND_181[6:0];
  _RAND_182 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfSrc1_p = _RAND_182[4:0];
  _RAND_183 = {1{`RANDOM}};
  toggle_9552_valid_reg = _RAND_183[4:0];
  _RAND_184 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfSrc2_p = _RAND_184[4:0];
  _RAND_185 = {1{`RANDOM}};
  toggle_9557_valid_reg = _RAND_185[4:0];
  _RAND_186 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfWen_p = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  toggle_9562_valid_reg = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  dataBuffer_1_ctrl_rfDest_p = _RAND_188[4:0];
  _RAND_189 = {1{`RANDOM}};
  toggle_9563_valid_reg = _RAND_189[4:0];
  _RAND_190 = {1{`RANDOM}};
  dataBuffer_1_ctrl_isNutCoreTrap_p = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  toggle_9568_valid_reg = _RAND_191[0:0];
  _RAND_192 = {2{`RANDOM}};
  dataBuffer_1_data_imm_p = _RAND_192[63:0];
  _RAND_193 = {2{`RANDOM}};
  toggle_9569_valid_reg = _RAND_193[63:0];
  _RAND_194 = {2{`RANDOM}};
  dataBuffer_2_cf_instr_p = _RAND_194[63:0];
  _RAND_195 = {2{`RANDOM}};
  toggle_9633_valid_reg = _RAND_195[63:0];
  _RAND_196 = {2{`RANDOM}};
  dataBuffer_2_cf_pc_p = _RAND_196[38:0];
  _RAND_197 = {2{`RANDOM}};
  toggle_9697_valid_reg = _RAND_197[38:0];
  _RAND_198 = {2{`RANDOM}};
  dataBuffer_2_cf_pnpc_p = _RAND_198[38:0];
  _RAND_199 = {2{`RANDOM}};
  toggle_9736_valid_reg = _RAND_199[38:0];
  _RAND_200 = {1{`RANDOM}};
  dataBuffer_2_cf_exceptionVec_1_p = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  toggle_9775_valid_reg = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  dataBuffer_2_cf_exceptionVec_2_p = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  toggle_9776_valid_reg = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  dataBuffer_2_cf_exceptionVec_12_p = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  toggle_9777_valid_reg = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_1_p = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  toggle_9778_valid_reg = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_3_p = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  toggle_9779_valid_reg = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_5_p = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  toggle_9780_valid_reg = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_7_p = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  toggle_9781_valid_reg = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_9_p = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  toggle_9782_valid_reg = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  dataBuffer_2_cf_intrVec_11_p = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  toggle_9783_valid_reg = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  dataBuffer_2_cf_brIdx_p = _RAND_218[3:0];
  _RAND_219 = {1{`RANDOM}};
  toggle_9784_valid_reg = _RAND_219[3:0];
  _RAND_220 = {1{`RANDOM}};
  dataBuffer_2_cf_crossBoundaryFault_p = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  toggle_9788_valid_reg = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  dataBuffer_2_ctrl_src1Type_p = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  toggle_9789_valid_reg = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  dataBuffer_2_ctrl_src2Type_p = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  toggle_9790_valid_reg = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  dataBuffer_2_ctrl_fuType_p = _RAND_226[2:0];
  _RAND_227 = {1{`RANDOM}};
  toggle_9791_valid_reg = _RAND_227[2:0];
  _RAND_228 = {1{`RANDOM}};
  dataBuffer_2_ctrl_fuOpType_p = _RAND_228[6:0];
  _RAND_229 = {1{`RANDOM}};
  toggle_9794_valid_reg = _RAND_229[6:0];
  _RAND_230 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfSrc1_p = _RAND_230[4:0];
  _RAND_231 = {1{`RANDOM}};
  toggle_9801_valid_reg = _RAND_231[4:0];
  _RAND_232 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfSrc2_p = _RAND_232[4:0];
  _RAND_233 = {1{`RANDOM}};
  toggle_9806_valid_reg = _RAND_233[4:0];
  _RAND_234 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfWen_p = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  toggle_9811_valid_reg = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  dataBuffer_2_ctrl_rfDest_p = _RAND_236[4:0];
  _RAND_237 = {1{`RANDOM}};
  toggle_9812_valid_reg = _RAND_237[4:0];
  _RAND_238 = {1{`RANDOM}};
  dataBuffer_2_ctrl_isNutCoreTrap_p = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  toggle_9817_valid_reg = _RAND_239[0:0];
  _RAND_240 = {2{`RANDOM}};
  dataBuffer_2_data_imm_p = _RAND_240[63:0];
  _RAND_241 = {2{`RANDOM}};
  toggle_9818_valid_reg = _RAND_241[63:0];
  _RAND_242 = {2{`RANDOM}};
  dataBuffer_3_cf_instr_p = _RAND_242[63:0];
  _RAND_243 = {2{`RANDOM}};
  toggle_9882_valid_reg = _RAND_243[63:0];
  _RAND_244 = {2{`RANDOM}};
  dataBuffer_3_cf_pc_p = _RAND_244[38:0];
  _RAND_245 = {2{`RANDOM}};
  toggle_9946_valid_reg = _RAND_245[38:0];
  _RAND_246 = {2{`RANDOM}};
  dataBuffer_3_cf_pnpc_p = _RAND_246[38:0];
  _RAND_247 = {2{`RANDOM}};
  toggle_9985_valid_reg = _RAND_247[38:0];
  _RAND_248 = {1{`RANDOM}};
  dataBuffer_3_cf_exceptionVec_1_p = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  toggle_10024_valid_reg = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  dataBuffer_3_cf_exceptionVec_2_p = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  toggle_10025_valid_reg = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  dataBuffer_3_cf_exceptionVec_12_p = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  toggle_10026_valid_reg = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_1_p = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  toggle_10027_valid_reg = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_3_p = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  toggle_10028_valid_reg = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_5_p = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  toggle_10029_valid_reg = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_7_p = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  toggle_10030_valid_reg = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_9_p = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  toggle_10031_valid_reg = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  dataBuffer_3_cf_intrVec_11_p = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  toggle_10032_valid_reg = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  dataBuffer_3_cf_brIdx_p = _RAND_266[3:0];
  _RAND_267 = {1{`RANDOM}};
  toggle_10033_valid_reg = _RAND_267[3:0];
  _RAND_268 = {1{`RANDOM}};
  dataBuffer_3_cf_crossBoundaryFault_p = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  toggle_10037_valid_reg = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  dataBuffer_3_ctrl_src1Type_p = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  toggle_10038_valid_reg = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  dataBuffer_3_ctrl_src2Type_p = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  toggle_10039_valid_reg = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  dataBuffer_3_ctrl_fuType_p = _RAND_274[2:0];
  _RAND_275 = {1{`RANDOM}};
  toggle_10040_valid_reg = _RAND_275[2:0];
  _RAND_276 = {1{`RANDOM}};
  dataBuffer_3_ctrl_fuOpType_p = _RAND_276[6:0];
  _RAND_277 = {1{`RANDOM}};
  toggle_10043_valid_reg = _RAND_277[6:0];
  _RAND_278 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfSrc1_p = _RAND_278[4:0];
  _RAND_279 = {1{`RANDOM}};
  toggle_10050_valid_reg = _RAND_279[4:0];
  _RAND_280 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfSrc2_p = _RAND_280[4:0];
  _RAND_281 = {1{`RANDOM}};
  toggle_10055_valid_reg = _RAND_281[4:0];
  _RAND_282 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfWen_p = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  toggle_10060_valid_reg = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  dataBuffer_3_ctrl_rfDest_p = _RAND_284[4:0];
  _RAND_285 = {1{`RANDOM}};
  toggle_10061_valid_reg = _RAND_285[4:0];
  _RAND_286 = {1{`RANDOM}};
  dataBuffer_3_ctrl_isNutCoreTrap_p = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  toggle_10066_valid_reg = _RAND_287[0:0];
  _RAND_288 = {2{`RANDOM}};
  dataBuffer_3_data_imm_p = _RAND_288[63:0];
  _RAND_289 = {2{`RANDOM}};
  toggle_10067_valid_reg = _RAND_289[63:0];
  _RAND_290 = {1{`RANDOM}};
  ringBufferHead_p = _RAND_290[1:0];
  _RAND_291 = {1{`RANDOM}};
  toggle_10131_valid_reg = _RAND_291[1:0];
  _RAND_292 = {1{`RANDOM}};
  ringBufferTail_p = _RAND_292[1:0];
  _RAND_293 = {1{`RANDOM}};
  toggle_10133_valid_reg = _RAND_293[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[5]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[6]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[7]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[8]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[9]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[10]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[11]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[12]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[13]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[14]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[15]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[16]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[17]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[18]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[19]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[20]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[21]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[22]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[23]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[24]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[25]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[26]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[27]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[28]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[29]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[30]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[31]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[32]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[33]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[34]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[35]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[36]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[37]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[38]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[39]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[40]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[41]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[42]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[43]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[44]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[45]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[46]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[47]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[48]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[49]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[50]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[51]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[52]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[53]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[54]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[55]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[56]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[57]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[58]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[59]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[60]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[61]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[62]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_instr_t[63]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[5]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[6]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[7]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[8]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[9]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[10]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[11]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[12]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[13]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[14]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[15]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[16]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[17]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[18]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[19]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[20]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[21]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[22]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[23]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[24]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[25]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[26]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[27]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[28]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[29]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[30]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[31]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[32]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[33]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[34]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[35]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[36]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[37]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pc_t[38]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[5]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[6]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[7]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[8]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[9]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[10]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[11]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[12]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[13]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[14]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[15]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[16]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[17]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[18]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[19]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[20]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[21]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[22]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[23]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[24]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[25]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[26]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[27]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[28]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[29]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[30]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[31]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[32]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[33]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[34]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[35]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[36]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[37]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_pnpc_t[38]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_exceptionVec_1_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_exceptionVec_2_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_exceptionVec_12_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_intrVec_1_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_intrVec_3_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_intrVec_5_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_intrVec_7_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_intrVec_9_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_intrVec_11_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_brIdx_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_brIdx_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_brIdx_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_brIdx_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_cf_crossBoundaryFault_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_src1Type_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_src2Type_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_fuType_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_fuType_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_fuType_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_fuOpType_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_fuOpType_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_fuOpType_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_fuOpType_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_fuOpType_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_fuOpType_t[5]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_fuOpType_t[6]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_rfSrc1_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_rfSrc1_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_rfSrc1_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_rfSrc1_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_rfSrc1_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_rfSrc2_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_rfSrc2_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_rfSrc2_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_rfSrc2_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_rfSrc2_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_rfWen_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_rfDest_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_rfDest_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_rfDest_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_rfDest_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_rfDest_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_ctrl_isNutCoreTrap_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[5]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[6]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[7]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[8]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[9]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[10]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[11]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[12]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[13]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[14]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[15]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[16]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[17]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[18]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[19]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[20]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[21]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[22]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[23]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[24]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[25]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[26]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[27]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[28]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[29]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[30]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[31]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[32]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[33]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[34]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[35]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[36]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[37]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[38]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[39]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[40]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[41]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[42]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[43]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[44]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[45]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[46]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[47]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[48]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[49]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[50]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[51]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[52]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[53]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[54]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[55]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[56]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[57]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[58]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[59]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[60]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[61]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[62]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_0_data_imm_t[63]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[5]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[6]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[7]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[8]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[9]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[10]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[11]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[12]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[13]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[14]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[15]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[16]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[17]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[18]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[19]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[20]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[21]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[22]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[23]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[24]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[25]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[26]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[27]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[28]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[29]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[30]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[31]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[32]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[33]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[34]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[35]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[36]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[37]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[38]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[39]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[40]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[41]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[42]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[43]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[44]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[45]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[46]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[47]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[48]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[49]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[50]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[51]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[52]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[53]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[54]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[55]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[56]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[57]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[58]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[59]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[60]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[61]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[62]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_instr_t[63]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[5]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[6]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[7]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[8]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[9]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[10]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[11]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[12]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[13]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[14]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[15]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[16]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[17]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[18]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[19]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[20]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[21]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[22]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[23]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[24]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[25]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[26]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[27]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[28]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[29]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[30]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[31]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[32]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[33]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[34]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[35]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[36]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[37]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pc_t[38]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[5]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[6]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[7]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[8]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[9]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[10]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[11]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[12]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[13]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[14]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[15]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[16]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[17]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[18]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[19]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[20]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[21]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[22]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[23]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[24]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[25]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[26]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[27]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[28]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[29]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[30]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[31]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[32]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[33]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[34]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[35]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[36]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[37]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_pnpc_t[38]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_exceptionVec_1_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_exceptionVec_2_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_exceptionVec_12_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_intrVec_1_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_intrVec_3_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_intrVec_5_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_intrVec_7_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_intrVec_9_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_intrVec_11_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_brIdx_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_brIdx_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_brIdx_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_brIdx_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_cf_crossBoundaryFault_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_src1Type_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_src2Type_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_fuType_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_fuType_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_fuType_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_fuOpType_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_fuOpType_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_fuOpType_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_fuOpType_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_fuOpType_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_fuOpType_t[5]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_fuOpType_t[6]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_rfSrc1_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_rfSrc1_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_rfSrc1_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_rfSrc1_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_rfSrc1_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_rfSrc2_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_rfSrc2_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_rfSrc2_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_rfSrc2_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_rfSrc2_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_rfWen_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_rfDest_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_rfDest_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_rfDest_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_rfDest_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_rfDest_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_ctrl_isNutCoreTrap_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[5]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[6]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[7]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[8]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[9]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[10]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[11]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[12]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[13]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[14]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[15]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[16]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[17]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[18]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[19]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[20]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[21]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[22]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[23]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[24]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[25]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[26]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[27]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[28]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[29]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[30]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[31]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[32]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[33]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[34]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[35]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[36]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[37]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[38]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[39]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[40]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[41]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[42]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[43]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[44]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[45]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[46]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[47]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[48]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[49]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[50]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[51]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[52]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[53]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[54]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[55]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[56]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[57]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[58]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[59]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[60]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[61]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[62]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_1_data_imm_t[63]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[5]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[6]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[7]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[8]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[9]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[10]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[11]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[12]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[13]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[14]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[15]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[16]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[17]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[18]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[19]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[20]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[21]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[22]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[23]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[24]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[25]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[26]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[27]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[28]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[29]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[30]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[31]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[32]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[33]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[34]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[35]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[36]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[37]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[38]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[39]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[40]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[41]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[42]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[43]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[44]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[45]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[46]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[47]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[48]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[49]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[50]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[51]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[52]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[53]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[54]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[55]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[56]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[57]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[58]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[59]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[60]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[61]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[62]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_instr_t[63]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[5]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[6]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[7]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[8]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[9]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[10]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[11]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[12]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[13]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[14]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[15]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[16]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[17]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[18]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[19]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[20]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[21]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[22]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[23]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[24]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[25]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[26]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[27]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[28]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[29]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[30]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[31]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[32]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[33]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[34]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[35]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[36]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[37]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pc_t[38]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[5]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[6]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[7]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[8]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[9]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[10]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[11]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[12]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[13]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[14]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[15]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[16]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[17]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[18]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[19]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[20]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[21]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[22]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[23]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[24]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[25]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[26]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[27]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[28]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[29]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[30]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[31]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[32]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[33]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[34]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[35]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[36]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[37]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_pnpc_t[38]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_exceptionVec_1_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_exceptionVec_2_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_exceptionVec_12_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_intrVec_1_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_intrVec_3_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_intrVec_5_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_intrVec_7_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_intrVec_9_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_intrVec_11_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_brIdx_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_brIdx_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_brIdx_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_brIdx_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_cf_crossBoundaryFault_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_src1Type_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_src2Type_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_fuType_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_fuType_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_fuType_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_fuOpType_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_fuOpType_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_fuOpType_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_fuOpType_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_fuOpType_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_fuOpType_t[5]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_fuOpType_t[6]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_rfSrc1_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_rfSrc1_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_rfSrc1_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_rfSrc1_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_rfSrc1_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_rfSrc2_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_rfSrc2_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_rfSrc2_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_rfSrc2_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_rfSrc2_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_rfWen_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_rfDest_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_rfDest_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_rfDest_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_rfDest_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_rfDest_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_ctrl_isNutCoreTrap_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[5]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[6]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[7]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[8]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[9]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[10]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[11]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[12]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[13]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[14]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[15]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[16]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[17]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[18]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[19]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[20]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[21]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[22]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[23]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[24]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[25]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[26]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[27]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[28]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[29]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[30]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[31]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[32]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[33]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[34]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[35]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[36]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[37]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[38]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[39]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[40]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[41]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[42]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[43]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[44]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[45]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[46]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[47]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[48]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[49]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[50]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[51]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[52]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[53]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[54]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[55]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[56]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[57]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[58]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[59]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[60]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[61]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[62]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_2_data_imm_t[63]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[5]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[6]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[7]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[8]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[9]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[10]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[11]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[12]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[13]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[14]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[15]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[16]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[17]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[18]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[19]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[20]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[21]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[22]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[23]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[24]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[25]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[26]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[27]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[28]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[29]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[30]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[31]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[32]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[33]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[34]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[35]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[36]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[37]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[38]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[39]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[40]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[41]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[42]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[43]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[44]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[45]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[46]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[47]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[48]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[49]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[50]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[51]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[52]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[53]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[54]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[55]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[56]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[57]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[58]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[59]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[60]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[61]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[62]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_instr_t[63]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[5]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[6]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[7]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[8]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[9]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[10]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[11]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[12]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[13]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[14]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[15]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[16]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[17]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[18]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[19]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[20]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[21]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[22]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[23]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[24]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[25]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[26]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[27]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[28]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[29]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[30]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[31]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[32]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[33]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[34]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[35]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[36]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[37]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pc_t[38]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[5]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[6]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[7]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[8]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[9]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[10]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[11]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[12]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[13]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[14]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[15]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[16]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[17]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[18]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[19]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[20]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[21]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[22]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[23]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[24]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[25]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[26]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[27]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[28]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[29]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[30]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[31]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[32]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[33]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[34]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[35]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[36]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[37]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_pnpc_t[38]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_exceptionVec_1_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_exceptionVec_2_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_exceptionVec_12_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_intrVec_1_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_intrVec_3_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_intrVec_5_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_intrVec_7_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_intrVec_9_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_intrVec_11_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_brIdx_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_brIdx_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_brIdx_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_brIdx_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_cf_crossBoundaryFault_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_src1Type_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_src2Type_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_fuType_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_fuType_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_fuType_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_fuOpType_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_fuOpType_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_fuOpType_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_fuOpType_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_fuOpType_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_fuOpType_t[5]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_fuOpType_t[6]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_rfSrc1_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_rfSrc1_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_rfSrc1_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_rfSrc1_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_rfSrc1_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_rfSrc2_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_rfSrc2_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_rfSrc2_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_rfSrc2_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_rfSrc2_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_rfWen_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_rfDest_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_rfDest_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_rfDest_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_rfDest_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_rfDest_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_ctrl_isNutCoreTrap_t); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[0]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[1]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[2]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[3]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[4]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[5]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[6]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[7]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[8]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[9]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[10]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[11]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[12]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[13]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[14]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[15]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[16]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[17]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[18]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[19]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[20]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[21]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[22]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[23]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[24]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[25]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[26]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[27]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[28]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[29]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[30]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[31]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[32]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[33]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[34]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[35]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[36]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[37]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[38]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[39]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[40]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[41]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[42]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[43]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[44]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[45]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[46]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[47]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[48]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[49]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[50]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[51]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[52]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[53]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[54]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[55]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[56]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[57]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[58]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[59]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[60]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[61]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[62]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(dataBuffer_3_data_imm_t[63]); // @[src/main/scala/utils/PipelineVector.scala 29:29]
    end
    //
    if (enToggle_past) begin
      cover(ringBufferHead_t[0]); // @[src/main/scala/utils/PipelineVector.scala 30:33]
    end
    //
    if (enToggle_past) begin
      cover(ringBufferHead_t[1]); // @[src/main/scala/utils/PipelineVector.scala 30:33]
    end
    //
    if (enToggle_past) begin
      cover(ringBufferTail_t[0]); // @[src/main/scala/utils/PipelineVector.scala 31:33]
    end
    //
    if (enToggle_past) begin
      cover(ringBufferTail_t[1]); // @[src/main/scala/utils/PipelineVector.scala 31:33]
    end
  end
endmodule
module CoherenceManager(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/system/Coherence.scala 31:14]
  input         io_in_req_valid, // @[src/main/scala/system/Coherence.scala 31:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/system/Coherence.scala 31:14]
  output        io_in_resp_valid, // @[src/main/scala/system/Coherence.scala 31:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/system/Coherence.scala 31:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/system/Coherence.scala 31:14]
  input         io_out_mem_req_ready, // @[src/main/scala/system/Coherence.scala 31:14]
  output        io_out_mem_req_valid, // @[src/main/scala/system/Coherence.scala 31:14]
  output [31:0] io_out_mem_req_bits_addr, // @[src/main/scala/system/Coherence.scala 31:14]
  output        io_out_mem_resp_ready, // @[src/main/scala/system/Coherence.scala 31:14]
  input         io_out_mem_resp_valid, // @[src/main/scala/system/Coherence.scala 31:14]
  input  [3:0]  io_out_mem_resp_bits_cmd, // @[src/main/scala/system/Coherence.scala 31:14]
  input  [63:0] io_out_mem_resp_bits_rdata // @[src/main/scala/system/Coherence.scala 31:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[src/main/scala/system/Coherence.scala 45:22]
  wire  inflight = state != 3'h0; // @[src/main/scala/system/Coherence.scala 46:24]
  wire  _reqLatch_T = ~inflight; // @[src/main/scala/system/Coherence.scala 52:42]
  reg [31:0] reqLatch_addr; // @[src/main/scala/system/Coherence.scala 52:27]
  wire  _io_out_mem_req_valid_T_1 = io_in_req_valid & _reqLatch_T; // @[src/main/scala/system/Coherence.scala 65:43]
  wire  _T_20 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_31 = io_in_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:26]
  wire [2:0] _GEN_14 = io_in_resp_valid & _T_31 ? 3'h0 : state; // @[src/main/scala/system/Coherence.scala 45:22 89:{60,68}]
  wire  _T_34 = io_out_mem_req_ready & io_out_mem_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _GEN_15 = _T_34 ? 3'h4 : state; // @[src/main/scala/system/Coherence.scala 45:22 94:{36,44}]
  wire  _T_36 = io_out_mem_resp_ready & io_out_mem_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_37 = io_out_mem_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:26]
  wire [2:0] _GEN_16 = _T_36 & _T_37 ? 3'h0 : state; // @[src/main/scala/system/Coherence.scala 96:101 45:22 96:93]
  wire [2:0] _GEN_17 = _T_36 ? 3'h0 : state; // @[src/main/scala/system/Coherence.scala 45:22 97:{57,65}]
  wire [2:0] _GEN_18 = 3'h5 == state ? _GEN_17 : state; // @[src/main/scala/system/Coherence.scala 74:18 45:22]
  wire [2:0] _GEN_19 = 3'h4 == state ? _GEN_16 : _GEN_18; // @[src/main/scala/system/Coherence.scala 74:18]
  wire [31:0] _GEN_20 = 3'h3 == state ? reqLatch_addr : io_in_req_bits_addr; // @[src/main/scala/system/Coherence.scala 74:18 59:23 92:27]
  wire  _GEN_25 = 3'h3 == state | _io_out_mem_req_valid_T_1; // @[src/main/scala/system/Coherence.scala 74:18 93:28]
  wire [2:0] _GEN_26 = 3'h3 == state ? _GEN_15 : _GEN_19; // @[src/main/scala/system/Coherence.scala 74:18]
  wire  _GEN_28 = 3'h2 == state ? 1'h0 : io_out_mem_resp_valid; // @[src/main/scala/system/Coherence.scala 72:14 74:18 88:16]
  wire [3:0] _GEN_29 = 3'h2 == state ? 4'h0 : io_out_mem_resp_bits_cmd; // @[src/main/scala/system/Coherence.scala 72:14 74:18 88:16]
  wire [63:0] _GEN_30 = 3'h2 == state ? 64'h0 : io_out_mem_resp_bits_rdata; // @[src/main/scala/system/Coherence.scala 72:14 74:18 88:16]
  wire [31:0] _GEN_32 = 3'h2 == state ? io_in_req_bits_addr : _GEN_20; // @[src/main/scala/system/Coherence.scala 74:18 59:23]
  wire  _GEN_37 = 3'h2 == state ? _io_out_mem_req_valid_T_1 : _GEN_25; // @[src/main/scala/system/Coherence.scala 74:18]
  wire  _GEN_40 = 3'h1 == state ? io_out_mem_resp_valid : _GEN_28; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  wire [3:0] _GEN_41 = 3'h1 == state ? io_out_mem_resp_bits_cmd : _GEN_29; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  wire [63:0] _GEN_42 = 3'h1 == state ? io_out_mem_resp_bits_rdata : _GEN_30; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  wire [31:0] _GEN_43 = 3'h1 == state ? io_in_req_bits_addr : _GEN_32; // @[src/main/scala/system/Coherence.scala 74:18 59:23]
  wire  _GEN_48 = 3'h1 == state ? _io_out_mem_req_valid_T_1 : _GEN_37; // @[src/main/scala/system/Coherence.scala 74:18]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [2:0] state_p; // @[src/main/scala/system/Coherence.scala 45:22]
  wire [2:0] state_t = state ^ state_p; // @[src/main/scala/system/Coherence.scala 45:22]
  wire  toggle_10135_clock;
  wire  toggle_10135_reset;
  wire [2:0] toggle_10135_valid;
  reg [2:0] toggle_10135_valid_reg;
  reg [31:0] reqLatch_addr_p; // @[src/main/scala/system/Coherence.scala 52:27]
  wire [31:0] reqLatch_addr_t = reqLatch_addr ^ reqLatch_addr_p; // @[src/main/scala/system/Coherence.scala 52:27]
  wire  toggle_10138_clock;
  wire  toggle_10138_reset;
  wire [31:0] toggle_10138_valid;
  reg [31:0] toggle_10138_valid_reg;
  GEN_w3_toggle #(.COVER_INDEX(10135)) toggle_10135 (
    .clock(toggle_10135_clock),
    .reset(toggle_10135_reset),
    .valid(toggle_10135_valid)
  );
  GEN_w32_toggle #(.COVER_INDEX(10138)) toggle_10138 (
    .clock(toggle_10138_clock),
    .reset(toggle_10138_reset),
    .valid(toggle_10138_valid)
  );
  assign io_in_req_ready = io_out_mem_req_ready & _reqLatch_T; // @[src/main/scala/system/Coherence.scala 66:43]
  assign io_in_resp_valid = 3'h0 == state ? io_out_mem_resp_valid : _GEN_40; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  assign io_in_resp_bits_cmd = 3'h0 == state ? io_out_mem_resp_bits_cmd : _GEN_41; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  assign io_in_resp_bits_rdata = 3'h0 == state ? io_out_mem_resp_bits_rdata : _GEN_42; // @[src/main/scala/system/Coherence.scala 72:14 74:18]
  assign io_out_mem_req_valid = 3'h0 == state ? _io_out_mem_req_valid_T_1 : _GEN_48; // @[src/main/scala/system/Coherence.scala 74:18]
  assign io_out_mem_req_bits_addr = 3'h0 == state ? io_in_req_bits_addr : _GEN_43; // @[src/main/scala/system/Coherence.scala 74:18 59:23]
  assign io_out_mem_resp_ready = 1'h1; // @[src/main/scala/system/Coherence.scala 72:14]
  assign toggle_10135_clock = clock;
  assign toggle_10135_reset = reset;
  assign toggle_10135_valid = state ^ toggle_10135_valid_reg;
  assign toggle_10138_clock = clock;
  assign toggle_10138_reset = reset;
  assign toggle_10138_valid = reqLatch_addr ^ toggle_10138_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/system/Coherence.scala 45:22]
      state <= 3'h0; // @[src/main/scala/system/Coherence.scala 45:22]
    end else if (3'h0 == state) begin // @[src/main/scala/system/Coherence.scala 74:18]
      if (_T_20) begin // @[src/main/scala/system/Coherence.scala 76:29]
        state <= 3'h4;
      end
    end else if (!(3'h1 == state)) begin // @[src/main/scala/system/Coherence.scala 74:18]
      if (3'h2 == state) begin // @[src/main/scala/system/Coherence.scala 74:18]
        state <= _GEN_14;
      end else begin
        state <= _GEN_26;
      end
    end
    if (~inflight) begin // @[src/main/scala/system/Coherence.scala 52:27]
      reqLatch_addr <= io_in_req_bits_addr; // @[src/main/scala/system/Coherence.scala 52:27]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    state_p <= state; // @[src/main/scala/system/Coherence.scala 45:22]
    toggle_10135_valid_reg <= state;
    reqLatch_addr_p <= reqLatch_addr; // @[src/main/scala/system/Coherence.scala 52:27]
    toggle_10138_valid_reg <= reqLatch_addr;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  reqLatch_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  state_p = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  toggle_10135_valid_reg = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  reqLatch_addr_p = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  toggle_10138_valid_reg = _RAND_5[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(1'h1); // @[src/main/scala/system/Coherence.scala 49:9]
    end
    //
    if (enToggle_past) begin
      cover(state_t[0]); // @[src/main/scala/system/Coherence.scala 45:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[1]); // @[src/main/scala/system/Coherence.scala 45:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[2]); // @[src/main/scala/system/Coherence.scala 45:22]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[0]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[1]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[2]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[3]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[4]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[5]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[6]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[7]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[8]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[9]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[10]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[11]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[12]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[13]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[14]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[15]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[16]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[17]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[18]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[19]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[20]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[21]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[22]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[23]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[24]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[25]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[26]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[27]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[28]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[29]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[30]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
    //
    if (enToggle_past) begin
      cover(reqLatch_addr_t[31]); // @[src/main/scala/system/Coherence.scala 52:27]
    end
  end
endmodule
module LockingArbiter_2(
  input         clock,
  input         reset,
  output        io_in_0_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_0_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_0_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_in_1_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_in_1_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [31:0] io_in_1_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [2:0]  io_in_1_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [3:0]  io_in_1_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [7:0]  io_in_1_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input  [63:0] io_in_1_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  input         io_out_ready, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_out_valid, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [2:0]  io_out_bits_size, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [3:0]  io_out_bits_cmd, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [7:0]  io_out_bits_wmask, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output [63:0] io_out_bits_wdata, // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
  output        io_chosen // @[src/main/scala/chisel3/util/Arbiter.scala 52:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] lockCount_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg  lockIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
  wire  locked = lockCount_value != 3'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 61:34]
  wire  wantsLock = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[src/main/scala/bus/simplebus/Crossbar.scala 94:62]
  wire  _T = io_out_ready & io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [2:0] _value_T_1 = lockCount_value + 3'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  io_chosen_choice = io_in_0_valid ? 1'h0 : 1'h1; // @[src/main/scala/chisel3/util/Arbiter.scala 103:{26,35} 101:41]
  wire  _T_2 = ~io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 45:78]
  wire  _io_in_0_ready_T_1 = locked ? ~lockIdx : 1'h1; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  wire  _io_in_1_ready_T_1 = locked ? lockIdx : _T_2; // @[src/main/scala/chisel3/util/Arbiter.scala 71:22]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [2:0] lockCount_value_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [2:0] lockCount_value_t = lockCount_value ^ lockCount_value_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  toggle_10170_clock;
  wire  toggle_10170_reset;
  wire [2:0] toggle_10170_valid;
  reg [2:0] toggle_10170_valid_reg;
  reg  lockIdx_p; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
  wire  lockIdx_t = lockIdx ^ lockIdx_p; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
  wire  toggle_10173_clock;
  wire  toggle_10173_reset;
  wire  toggle_10173_valid;
  reg  toggle_10173_valid_reg;
  GEN_w3_toggle #(.COVER_INDEX(10170)) toggle_10170 (
    .clock(toggle_10170_clock),
    .reset(toggle_10170_reset),
    .valid(toggle_10170_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10173)) toggle_10173 (
    .clock(toggle_10173_clock),
    .reset(toggle_10173_reset),
    .valid(toggle_10173_valid)
  );
  assign io_in_0_ready = _io_in_0_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_in_1_ready = _io_in_1_ready_T_1 & io_out_ready; // @[src/main/scala/chisel3/util/Arbiter.scala 71:56]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[src/main/scala/chisel3/util/Arbiter.scala 55:{16,16}]
  assign io_out_bits_addr = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_size = io_chosen ? io_in_1_bits_size : 3'h3; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_cmd = io_chosen ? io_in_1_bits_cmd : 4'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wmask = io_chosen ? io_in_1_bits_wmask : 8'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_out_bits_wdata = io_chosen ? io_in_1_bits_wdata : 64'h0; // @[src/main/scala/chisel3/util/Arbiter.scala 56:{15,15}]
  assign io_chosen = locked ? lockIdx : io_chosen_choice; // @[src/main/scala/chisel3/util/Arbiter.scala 54:13 69:{18,30}]
  assign toggle_10170_clock = clock;
  assign toggle_10170_reset = reset;
  assign toggle_10170_valid = lockCount_value ^ toggle_10170_valid_reg;
  assign toggle_10173_clock = clock;
  assign toggle_10173_reset = reset;
  assign toggle_10173_valid = lockIdx ^ toggle_10173_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      lockCount_value <= 3'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockCount_value <= _value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (_T & wantsLock) begin // @[src/main/scala/chisel3/util/Arbiter.scala 64:36]
      lockIdx <= io_chosen; // @[src/main/scala/chisel3/util/Arbiter.scala 65:15]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    lockCount_value_p <= lockCount_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    toggle_10170_valid_reg <= lockCount_value;
    lockIdx_p <= lockIdx; // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
    toggle_10173_valid_reg <= lockIdx;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lockCount_value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  lockIdx = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  lockCount_value_p = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  toggle_10170_valid_reg = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  lockIdx_p = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  toggle_10173_valid_reg = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(lockCount_value_t[0]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(lockCount_value_t[1]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(lockCount_value_t[2]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(lockIdx_t); // @[src/main/scala/chisel3/util/Arbiter.scala 60:22]
    end
  end
endmodule
module SimpleBusCrossbarNto1_2(
  input         clock,
  input         reset,
  output        io_in_0_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_0_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_0_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_0_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_in_0_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_0_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_1_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_in_1_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [31:0] io_in_1_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [2:0]  io_in_1_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_in_1_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [7:0]  io_in_1_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_in_1_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_in_1_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_in_1_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_in_1_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_out_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_out_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [2:0]  io_out_req_bits_size, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  output        io_out_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input         io_out_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [3:0]  io_out_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
  input  [63:0] io_out_resp_bits_rdata // @[src/main/scala/bus/simplebus/Crossbar.scala 86:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_reset; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_0_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_in_1_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [2:0] inputArb_io_in_1_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_in_1_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_out_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_out_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [2:0] inputArb_io_out_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  wire  inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
  reg [1:0] state; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
  wire  _T_1 = ~inputArb_io_out_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:18]
  wire  _T_4 = ~inputArb_io_out_bits_cmd[0] & ~inputArb_io_out_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  reg  inflightSrc; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
  wire  _io_out_req_valid_T = state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 103:47]
  wire  _T_15 = inputArb_io_out_ready & inputArb_io_out_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_21 = inputArb_io_out_bits_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire  _T_22 = inputArb_io_out_bits_cmd == 4'h1; // @[src/main/scala/bus/simplebus/SimpleBus.scala 77:29]
  wire [1:0] _GEN_4 = _T_21 | _T_22 ? 2'h2 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 118:{80,88} 92:22]
  wire  _T_25 = io_out_resp_ready & io_out_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _T_26 = io_out_resp_bits_cmd == 4'h6; // @[src/main/scala/bus/simplebus/SimpleBus.scala 91:26]
  wire [1:0] _GEN_9 = _T_25 ? 2'h0 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 122:{50,58} 92:22]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [1:0] state_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
  wire [1:0] state_t = state ^ state_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
  wire  toggle_10174_clock;
  wire  toggle_10174_reset;
  wire [1:0] toggle_10174_valid;
  reg [1:0] toggle_10174_valid_reg;
  reg  inflightSrc_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
  wire  inflightSrc_t = inflightSrc ^ inflightSrc_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
  wire  toggle_10176_clock;
  wire  toggle_10176_reset;
  wire  toggle_10176_valid;
  reg  toggle_10176_valid_reg;
  LockingArbiter_2 inputArb ( // @[src/main/scala/bus/simplebus/Crossbar.scala 95:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_size(inputArb_io_in_1_bits_size),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(inputArb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_size(inputArb_io_out_bits_size),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  GEN_w2_toggle #(.COVER_INDEX(10174)) toggle_10174 (
    .clock(toggle_10174_clock),
    .reset(toggle_10174_reset),
    .valid(toggle_10174_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10176)) toggle_10176 (
    .clock(toggle_10176_clock),
    .reset(toggle_10176_reset),
    .valid(toggle_10176_valid)
  );
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_0_resp_valid = ~inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_0_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign io_in_1_resp_valid = inflightSrc & io_out_resp_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 109:{13,13} 107:26]
  assign io_in_1_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 106:25]
  assign io_out_req_valid = inputArb_io_out_valid & state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 103:37]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_size = inputArb_io_out_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 101:19]
  assign io_out_resp_ready = 1'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 110:{13,13}]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_size = io_in_1_req_bits_size; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_wmask = io_in_1_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 96:68]
  assign inputArb_io_out_ready = io_out_req_ready & _io_out_req_valid_T; // @[src/main/scala/bus/simplebus/Crossbar.scala 104:37]
  assign toggle_10174_clock = clock;
  assign toggle_10174_reset = reset;
  assign toggle_10174_valid = state ^ toggle_10174_valid_reg;
  assign toggle_10176_clock = clock;
  assign toggle_10176_reset = reset;
  assign toggle_10176_valid = inflightSrc ^ toggle_10176_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
      state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_15) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:29]
        if (_T_4) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 117:38]
          state <= 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 117:46]
        end else begin
          state <= _GEN_4;
        end
      end
    end else if (2'h1 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_25 & _T_26) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 121:82]
        state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 121:90]
      end
    end else if (2'h2 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      state <= _GEN_9;
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
      inflightSrc <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 113:18]
      if (_T_15) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 115:29]
        inflightSrc <= inputArb_io_chosen; // @[src/main/scala/bus/simplebus/Crossbar.scala 116:21]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(inputArb_io_out_valid & ~_T_4 & _T_1))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Crossbar.scala:98 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"
            ); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    state_p <= state; // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
    toggle_10174_valid_reg <= state;
    inflightSrc_p <= inflightSrc; // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
    toggle_10176_valid_reg <= inflightSrc;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  inflightSrc = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_p = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  toggle_10174_valid_reg = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  inflightSrc_p = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  toggle_10176_valid_reg = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~(inputArb_io_out_valid & ~_T_4 & _T_1)); // @[src/main/scala/bus/simplebus/Crossbar.scala 98:9]
    end
    //
    if (enToggle_past) begin
      cover(state_t[0]); // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[1]); // @[src/main/scala/bus/simplebus/Crossbar.scala 92:22]
    end
    //
    if (enToggle_past) begin
      cover(inflightSrc_t); // @[src/main/scala/bus/simplebus/Crossbar.scala 99:28]
    end
  end
endmodule
module AXI42SimpleBusConverter(
  input   clock,
  input   reset
);
endmodule
module SimpleBus2MemPortConverter(
  input   clock,
  input   reset
);
endmodule
module SimpleBusAddressMapper(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [2:0]  io_in_req_bits_size, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input         io_out_req_ready, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output        io_out_req_valid, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [31:0] io_out_req_bits_addr, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [2:0]  io_out_req_bits_size, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [3:0]  io_out_req_bits_cmd, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [7:0]  io_out_req_bits_wmask, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  output [63:0] io_out_req_bits_wdata, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input         io_out_resp_valid, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [3:0]  io_out_resp_bits_cmd, // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
  input  [63:0] io_out_resp_bits_rdata // @[src/main/scala/bus/simplebus/AddressMapper.scala 26:14]
);
  assign io_in_req_ready = io_out_req_ready; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_in_resp_valid = io_out_resp_valid; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_in_resp_bits_cmd = io_out_resp_bits_cmd; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_valid = io_in_req_valid; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_bits_size = io_in_req_bits_size; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
  assign io_out_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/AddressMapper.scala 31:10]
endmodule
module SimpleBus2AXI4Converter(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [2:0]  io_in_req_bits_size, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_aw_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_out_w_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_w_bits_strb, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_bits_last, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_ar_bits_len, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [2:0]  io_out_ar_bits_size, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_out_r_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_bits_last // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] _io_out_ar_bits_len_T_1 = io_in_req_bits_cmd[1] ? 3'h7 : 3'h0; // @[src/main/scala/bus/simplebus/ToAXI4.scala 169:30]
  wire  _io_out_w_bits_last_T = io_in_req_bits_cmd == 4'h7; // @[src/main/scala/bus/simplebus/SimpleBus.scala 78:27]
  wire  _io_out_w_bits_last_T_1 = io_in_req_bits_cmd == 4'h1; // @[src/main/scala/bus/simplebus/SimpleBus.scala 77:29]
  wire [2:0] _io_in_resp_bits_cmd_T = io_out_r_bits_last ? 3'h6 : 3'h0; // @[src/main/scala/bus/simplebus/ToAXI4.scala 184:28]
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 & io_out_w_bits_last | awAck & wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 189:53]
  wire  _wAck_T_1 = _wSend_T_1 & io_out_w_bits_last; // @[src/main/scala/bus/simplebus/ToAXI4.scala 188:41]
  wire  _GEN_2 = _wAck_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wen_T_1 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  _io_out_ar_valid_T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _io_out_aw_valid_T_1 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  wire  _io_out_w_valid_T_2 = ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:36]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  awAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  awAck_t = awAck ^ awAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10177_clock;
  wire  toggle_10177_reset;
  wire  toggle_10177_valid;
  reg  toggle_10177_valid_reg;
  reg  wAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wAck_t = wAck ^ wAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10178_clock;
  wire  toggle_10178_reset;
  wire  toggle_10178_valid;
  reg  toggle_10178_valid_reg;
  reg  wen_p; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  wen_t = wen ^ wen_p; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  toggle_10179_clock;
  wire  toggle_10179_reset;
  wire  toggle_10179_valid;
  reg  toggle_10179_valid_reg;
  GEN_w1_toggle #(.COVER_INDEX(10177)) toggle_10177 (
    .clock(toggle_10177_clock),
    .reset(toggle_10177_reset),
    .valid(toggle_10177_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10178)) toggle_10178 (
    .clock(toggle_10178_clock),
    .reset(toggle_10178_reset),
    .valid(toggle_10178_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10179)) toggle_10179 (
    .clock(toggle_10179_clock),
    .reset(toggle_10179_reset),
    .valid(toggle_10179_valid)
  );
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _io_out_w_valid_T_2 & io_out_w_ready : 1'h1; // @[src/main/scala/bus/simplebus/ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 199:25]
  assign io_in_resp_bits_cmd = {{1'd0}, _io_in_resp_bits_cmd_T}; // @[src/main/scala/bus/simplebus/ToAXI4.scala 184:22]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 183:23]
  assign io_out_aw_valid = _io_out_aw_valid_T_1 & ~awAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 193:33]
  assign io_out_aw_bits_addr = io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_w_valid = _io_out_aw_valid_T_1 & ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:33]
  assign io_out_w_bits_data = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 160:10]
  assign io_out_w_bits_strb = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 161:10]
  assign io_out_w_bits_last = _io_out_w_bits_last_T | _io_out_w_bits_last_T_1; // @[src/main/scala/bus/simplebus/ToAXI4.scala 177:54]
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 158:12]
  assign io_out_ar_bits_len = {{5'd0}, _io_out_ar_bits_len_T_1}; // @[src/main/scala/bus/simplebus/ToAXI4.scala 169:24]
  assign io_out_ar_bits_size = io_in_req_bits_size; // @[src/main/scala/bus/simplebus/ToAXI4.scala 170:24]
  assign toggle_10177_clock = clock;
  assign toggle_10177_reset = reset;
  assign toggle_10177_valid = awAck ^ toggle_10177_valid_reg;
  assign toggle_10178_clock = clock;
  assign toggle_10178_reset = reset;
  assign toggle_10178_valid = wAck ^ toggle_10178_valid_reg;
  assign toggle_10179_clock = clock;
  assign toggle_10179_reset = reset;
  assign toggle_10179_valid = wen ^ toggle_10179_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_2;
    end
    if (_wen_T_1) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
      wen <= io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    awAck_p <= awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10177_valid_reg <= awAck;
    wAck_p <= wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10178_valid_reg <= wAck;
    wen_p <= wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    toggle_10179_valid_reg <= wen;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  awAck_p = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  toggle_10177_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  wAck_p = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  toggle_10178_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  wen_p = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  toggle_10179_valid_reg = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(1'h1); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
    end
    //
    if (enToggle_past) begin
      cover(awAck_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(wAck_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(wen_t); // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
  end
endmodule
module SimpleBusCrossbar1toN(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_0_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_0_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_0_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_0_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_0_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_0_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_0_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_0_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_0_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_1_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_1_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_1_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_1_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_1_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_1_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_1_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_1_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_1_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_2_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_2_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_2_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_2_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_2_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_2_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_2_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_2_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [3:0]  io_out_2_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_2_resp_bits_rdata // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
  wire  outMatchVec_0 = io_in_req_bits_addr >= 32'h38000000 & io_in_req_bits_addr < 32'h38010000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_1 = io_in_req_bits_addr >= 32'h3c000000 & io_in_req_bits_addr < 32'h40000000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_2 = io_in_req_bits_addr >= 32'h40000000 & io_in_req_bits_addr < 32'h80000000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire [2:0] _outSelVec_enc_T = outMatchVec_2 ? 3'h4 : 3'h0; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _outSelVec_enc_T_1 = outMatchVec_1 ? 3'h2 : _outSelVec_enc_T; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] outSelVec_enc = outMatchVec_0 ? 3'h1 : _outSelVec_enc_T_1; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire  outSelVec_0 = outSelVec_enc[0]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_1 = outSelVec_enc[1]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_2 = outSelVec_enc[2]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  _outSelRespVec_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _outSelRespVec_T_1 = state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 41:59]
  wire  _outSelRespVec_T_2 = _outSelRespVec_T & state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 41:50]
  reg  outSelRespVec_0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_2; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire [2:0] _reqInvalidAddr_T = {outSelVec_2,outSelVec_1,outSelVec_0}; // @[src/main/scala/bus/simplebus/Crossbar.scala 42:54]
  wire  reqInvalidAddr = io_in_req_valid & ~(|_reqInvalidAddr_T); // @[src/main/scala/bus/simplebus/Crossbar.scala 42:40]
  wire [1:0] _GEN_5 = io_in_resp_valid ? 2'h0 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22 56:{44,52}]
  wire  _io_in_req_ready_T_4 = outSelVec_0 & io_out_0_req_ready | outSelVec_1 & io_out_1_req_ready | outSelVec_2 &
    io_out_2_req_ready; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_in_resp_valid_T_4 = outSelRespVec_0 & io_out_0_resp_valid | outSelRespVec_1 & io_out_1_resp_valid |
    outSelRespVec_2 & io_out_2_resp_valid; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T = outSelRespVec_0 ? io_out_0_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_1 = outSelRespVec_1 ? io_out_1_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_2 = outSelRespVec_2 ? io_out_2_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_3 = _io_in_resp_bits_T | _io_in_resp_bits_T_1; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_5 = outSelRespVec_0 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_6 = outSelRespVec_1 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_7 = outSelRespVec_2 ? io_out_2_resp_bits_cmd : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_8 = _io_in_resp_bits_T_5 | _io_in_resp_bits_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [1:0] state_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
  wire [1:0] state_t = state ^ state_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
  wire  toggle_10180_clock;
  wire  toggle_10180_reset;
  wire [1:0] toggle_10180_valid;
  reg [1:0] toggle_10180_valid_reg;
  reg  outSelRespVec_0_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire  outSelRespVec_0_t = outSelRespVec_0 ^ outSelRespVec_0_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire  toggle_10182_clock;
  wire  toggle_10182_reset;
  wire  toggle_10182_valid;
  reg  toggle_10182_valid_reg;
  reg  outSelRespVec_1_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire  outSelRespVec_1_t = outSelRespVec_1 ^ outSelRespVec_1_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire  toggle_10183_clock;
  wire  toggle_10183_reset;
  wire  toggle_10183_valid;
  reg  toggle_10183_valid_reg;
  reg  outSelRespVec_2_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire  outSelRespVec_2_t = outSelRespVec_2 ^ outSelRespVec_2_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire  toggle_10184_clock;
  wire  toggle_10184_reset;
  wire  toggle_10184_valid;
  reg  toggle_10184_valid_reg;
  GEN_w2_toggle #(.COVER_INDEX(10180)) toggle_10180 (
    .clock(toggle_10180_clock),
    .reset(toggle_10180_reset),
    .valid(toggle_10180_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10182)) toggle_10182 (
    .clock(toggle_10182_clock),
    .reset(toggle_10182_reset),
    .valid(toggle_10182_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10183)) toggle_10183 (
    .clock(toggle_10183_clock),
    .reset(toggle_10183_reset),
    .valid(toggle_10183_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10184)) toggle_10184 (
    .clock(toggle_10184_clock),
    .reset(toggle_10184_reset),
    .valid(toggle_10184_valid)
  );
  assign io_in_req_ready = _io_in_req_ready_T_4 | reqInvalidAddr; // @[src/main/scala/bus/simplebus/Crossbar.scala 61:64]
  assign io_in_resp_valid = _io_in_resp_valid_T_4 | state == 2'h2; // @[src/main/scala/bus/simplebus/Crossbar.scala 71:70]
  assign io_in_resp_bits_cmd = _io_in_resp_bits_T_8 | _io_in_resp_bits_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_in_resp_bits_rdata = _io_in_resp_bits_T_3 | _io_in_resp_bits_T_2; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_0_req_valid = outSelVec_0 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_0_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_resp_ready = outSelRespVec_0 & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_1_req_valid = outSelVec_1 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_1_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_resp_ready = outSelRespVec_1 & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_2_req_valid = outSelVec_2 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_2_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_resp_ready = outSelRespVec_2 & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign toggle_10180_clock = clock;
  assign toggle_10180_reset = reset;
  assign toggle_10180_valid = state ^ toggle_10180_valid_reg;
  assign toggle_10182_clock = clock;
  assign toggle_10182_reset = reset;
  assign toggle_10182_valid = outSelRespVec_0 ^ toggle_10182_valid_reg;
  assign toggle_10183_clock = clock;
  assign toggle_10183_reset = reset;
  assign toggle_10183_valid = outSelRespVec_1 ^ toggle_10183_valid_reg;
  assign toggle_10184_clock = clock;
  assign toggle_10184_reset = reset;
  assign toggle_10184_valid = outSelRespVec_2 ^ toggle_10184_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
      state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      if (reqInvalidAddr) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 54:29]
        state <= 2'h2; // @[src/main/scala/bus/simplebus/Crossbar.scala 54:37]
      end else if (_outSelRespVec_T) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 53:31]
        state <= 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 53:39]
      end
    end else if (2'h1 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      state <= _GEN_5;
    end else if (2'h2 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      state <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_0 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_0 <= outSelVec_0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_1 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_1 <= outSelVec_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_2 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_2 <= outSelVec_2; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~reqInvalidAddr)) begin
          $fwrite(32'h80000002,
            "Assertion failed: address decode error, bad addr = 0x%x\n\n    at Crossbar.scala:49 assert(!reqInvalidAddr, \"address decode error, bad addr = 0x%%%%x\\n\", addr)\n"
            ,io_in_req_bits_addr); // @[src/main/scala/bus/simplebus/Crossbar.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    state_p <= state; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
    toggle_10180_valid_reg <= state;
    outSelRespVec_0_p <= outSelRespVec_0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    toggle_10182_valid_reg <= outSelRespVec_0;
    outSelRespVec_1_p <= outSelRespVec_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    toggle_10183_valid_reg <= outSelRespVec_1;
    outSelRespVec_2_p <= outSelRespVec_2; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    toggle_10184_valid_reg <= outSelRespVec_2;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  outSelRespVec_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  outSelRespVec_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  outSelRespVec_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state_p = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  toggle_10180_valid_reg = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  outSelRespVec_0_p = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  toggle_10182_valid_reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  outSelRespVec_1_p = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  toggle_10183_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  outSelRespVec_2_p = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  toggle_10184_valid_reg = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~reqInvalidAddr); // @[src/main/scala/bus/simplebus/Crossbar.scala 49:9]
    end
    //
    if (enToggle_past) begin
      cover(state_t[0]); // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[1]); // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(outSelRespVec_0_t); // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    //
    if (enToggle_past) begin
      cover(outSelRespVec_1_t); // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    //
    if (enToggle_past) begin
      cover(outSelRespVec_2_t); // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
  end
endmodule
module AXI4CLINT(
  input         clock,
  input         reset,
  output        io__in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io__in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io__in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io__in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io__in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io__in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__extra_mtip, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__extra_msip, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         isWFI_0,
  output        io_extra_mtip,
  output        io_extra_msip
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] _fullMask_T_8 = io__in_w_bits_strb[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_9 = io__in_w_bits_strb[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_10 = io__in_w_bits_strb[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_11 = io__in_w_bits_strb[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_12 = io__in_w_bits_strb[4] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_13 = io__in_w_bits_strb[5] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_14 = io__in_w_bits_strb[6] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_15 = io__in_w_bits_strb[7] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [63:0] fullMask = {_fullMask_T_15,_fullMask_T_14,_fullMask_T_13,_fullMask_T_12,_fullMask_T_11,_fullMask_T_10,
    _fullMask_T_9,_fullMask_T_8}; // @[src/main/scala/utils/BitUtils.scala 27:27]
  wire  _r_busy_T = io__in_ar_ready & io__in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _r_busy_T_1 = io__in_r_ready & io__in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _r_busy_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_2 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io__in_aw_ready & io__in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io__in_b_ready & io__in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _w_busy_T | _GEN_4; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io__in_w_ready & io__in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [63:0] mtime; // @[src/main/scala/device/AXI4CLINT.scala 32:22]
  reg [63:0] mtimecmp; // @[src/main/scala/device/AXI4CLINT.scala 33:25]
  reg [63:0] msip; // @[src/main/scala/device/AXI4CLINT.scala 34:21]
  reg [63:0] freq_reg; // @[src/main/scala/device/AXI4CLINT.scala 37:25]
  wire [15:0] freq = freq_reg[15:0]; // @[src/main/scala/device/AXI4CLINT.scala 38:22]
  reg [63:0] inc_reg; // @[src/main/scala/device/AXI4CLINT.scala 39:24]
  wire [15:0] inc = inc_reg[15:0]; // @[src/main/scala/device/AXI4CLINT.scala 40:20]
  reg [15:0] cnt; // @[src/main/scala/device/AXI4CLINT.scala 42:20]
  wire [15:0] nextCnt = cnt + 16'h1; // @[src/main/scala/device/AXI4CLINT.scala 43:21]
  wire  tick = nextCnt == freq; // @[src/main/scala/device/AXI4CLINT.scala 45:23]
  wire [63:0] _GEN_28 = {{48'd0}, inc}; // @[src/main/scala/device/AXI4CLINT.scala 46:32]
  wire [63:0] _mtime_T_1 = mtime + _GEN_28; // @[src/main/scala/device/AXI4CLINT.scala 46:32]
  wire [63:0] _mtime_T_3 = mtime + 64'h186a0; // @[src/main/scala/device/AXI4CLINT.scala 51:35]
  wire  _io_in_r_bits_data_T = 16'h0 == io__in_ar_bits_addr[15:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_1 = 16'h8000 == io__in_ar_bits_addr[15:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_2 = 16'hbff8 == io__in_ar_bits_addr[15:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_3 = 16'h8008 == io__in_ar_bits_addr[15:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_4 = 16'h4000 == io__in_ar_bits_addr[15:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [63:0] _io_in_r_bits_data_T_5 = _io_in_r_bits_data_T ? msip : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_6 = _io_in_r_bits_data_T_1 ? freq_reg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_7 = _io_in_r_bits_data_T_2 ? mtime : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_8 = _io_in_r_bits_data_T_3 ? inc_reg : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_9 = _io_in_r_bits_data_T_4 ? mtimecmp : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_10 = _io_in_r_bits_data_T_5 | _io_in_r_bits_data_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_11 = _io_in_r_bits_data_T_10 | _io_in_r_bits_data_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_r_bits_data_T_12 = _io_in_r_bits_data_T_11 | _io_in_r_bits_data_T_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _msip_T = io__in_w_bits_data & fullMask; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [63:0] _msip_T_1 = ~fullMask; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [63:0] _msip_T_2 = msip & _msip_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _msip_T_3 = _msip_T | _msip_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _freq_reg_T_2 = freq_reg & _msip_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _freq_reg_T_3 = _msip_T | _freq_reg_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _mtime_T_6 = mtime & _msip_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mtime_T_7 = _msip_T | _mtime_T_6; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _inc_reg_T_2 = inc_reg & _msip_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _inc_reg_T_3 = _msip_T | _inc_reg_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] _mtimecmp_T_2 = mtimecmp & _msip_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [63:0] _mtimecmp_T_3 = _msip_T | _mtimecmp_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  reg  io_extra_mtip_REG; // @[src/main/scala/device/AXI4CLINT.scala 66:31]
  reg  io_extra_msip_REG; // @[src/main/scala/device/AXI4CLINT.scala 67:31]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  r_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  r_busy_t = r_busy ^ r_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10185_clock;
  wire  toggle_10185_reset;
  wire  toggle_10185_valid;
  reg  toggle_10185_valid_reg;
  reg  ren_REG_p; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  ren_REG_t = ren_REG ^ ren_REG_p; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  toggle_10186_clock;
  wire  toggle_10186_reset;
  wire  toggle_10186_valid;
  reg  toggle_10186_valid_reg;
  reg  io_in_r_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  io_in_r_valid_r_t = io_in_r_valid_r ^ io_in_r_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10187_clock;
  wire  toggle_10187_reset;
  wire  toggle_10187_valid;
  reg  toggle_10187_valid_reg;
  reg  w_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  w_busy_t = w_busy ^ w_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10188_clock;
  wire  toggle_10188_reset;
  wire  toggle_10188_valid;
  reg  toggle_10188_valid_reg;
  reg  io_in_b_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  io_in_b_valid_r_t = io_in_b_valid_r ^ io_in_b_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10189_clock;
  wire  toggle_10189_reset;
  wire  toggle_10189_valid;
  reg  toggle_10189_valid_reg;
  reg [63:0] mtime_p; // @[src/main/scala/device/AXI4CLINT.scala 32:22]
  wire [63:0] mtime_t = mtime ^ mtime_p; // @[src/main/scala/device/AXI4CLINT.scala 32:22]
  wire  toggle_10190_clock;
  wire  toggle_10190_reset;
  wire [63:0] toggle_10190_valid;
  reg [63:0] toggle_10190_valid_reg;
  reg [63:0] mtimecmp_p; // @[src/main/scala/device/AXI4CLINT.scala 33:25]
  wire [63:0] mtimecmp_t = mtimecmp ^ mtimecmp_p; // @[src/main/scala/device/AXI4CLINT.scala 33:25]
  wire  toggle_10254_clock;
  wire  toggle_10254_reset;
  wire [63:0] toggle_10254_valid;
  reg [63:0] toggle_10254_valid_reg;
  reg [63:0] msip_p; // @[src/main/scala/device/AXI4CLINT.scala 34:21]
  wire [63:0] msip_t = msip ^ msip_p; // @[src/main/scala/device/AXI4CLINT.scala 34:21]
  wire  toggle_10318_clock;
  wire  toggle_10318_reset;
  wire [63:0] toggle_10318_valid;
  reg [63:0] toggle_10318_valid_reg;
  reg [63:0] freq_reg_p; // @[src/main/scala/device/AXI4CLINT.scala 37:25]
  wire [63:0] freq_reg_t = freq_reg ^ freq_reg_p; // @[src/main/scala/device/AXI4CLINT.scala 37:25]
  wire  toggle_10382_clock;
  wire  toggle_10382_reset;
  wire [63:0] toggle_10382_valid;
  reg [63:0] toggle_10382_valid_reg;
  reg [63:0] inc_reg_p; // @[src/main/scala/device/AXI4CLINT.scala 39:24]
  wire [63:0] inc_reg_t = inc_reg ^ inc_reg_p; // @[src/main/scala/device/AXI4CLINT.scala 39:24]
  wire  toggle_10446_clock;
  wire  toggle_10446_reset;
  wire [63:0] toggle_10446_valid;
  reg [63:0] toggle_10446_valid_reg;
  reg [15:0] cnt_p; // @[src/main/scala/device/AXI4CLINT.scala 42:20]
  wire [15:0] cnt_t = cnt ^ cnt_p; // @[src/main/scala/device/AXI4CLINT.scala 42:20]
  wire  toggle_10510_clock;
  wire  toggle_10510_reset;
  wire [15:0] toggle_10510_valid;
  reg [15:0] toggle_10510_valid_reg;
  reg  io_extra_mtip_REG_p; // @[src/main/scala/device/AXI4CLINT.scala 66:31]
  wire  io_extra_mtip_REG_t = io_extra_mtip_REG ^ io_extra_mtip_REG_p; // @[src/main/scala/device/AXI4CLINT.scala 66:31]
  wire  toggle_10526_clock;
  wire  toggle_10526_reset;
  wire  toggle_10526_valid;
  reg  toggle_10526_valid_reg;
  reg  io_extra_msip_REG_p; // @[src/main/scala/device/AXI4CLINT.scala 67:31]
  wire  io_extra_msip_REG_t = io_extra_msip_REG ^ io_extra_msip_REG_p; // @[src/main/scala/device/AXI4CLINT.scala 67:31]
  wire  toggle_10527_clock;
  wire  toggle_10527_reset;
  wire  toggle_10527_valid;
  reg  toggle_10527_valid_reg;
  GEN_w1_toggle #(.COVER_INDEX(10185)) toggle_10185 (
    .clock(toggle_10185_clock),
    .reset(toggle_10185_reset),
    .valid(toggle_10185_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10186)) toggle_10186 (
    .clock(toggle_10186_clock),
    .reset(toggle_10186_reset),
    .valid(toggle_10186_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10187)) toggle_10187 (
    .clock(toggle_10187_clock),
    .reset(toggle_10187_reset),
    .valid(toggle_10187_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10188)) toggle_10188 (
    .clock(toggle_10188_clock),
    .reset(toggle_10188_reset),
    .valid(toggle_10188_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10189)) toggle_10189 (
    .clock(toggle_10189_clock),
    .reset(toggle_10189_reset),
    .valid(toggle_10189_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(10190)) toggle_10190 (
    .clock(toggle_10190_clock),
    .reset(toggle_10190_reset),
    .valid(toggle_10190_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(10254)) toggle_10254 (
    .clock(toggle_10254_clock),
    .reset(toggle_10254_reset),
    .valid(toggle_10254_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(10318)) toggle_10318 (
    .clock(toggle_10318_clock),
    .reset(toggle_10318_reset),
    .valid(toggle_10318_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(10382)) toggle_10382 (
    .clock(toggle_10382_clock),
    .reset(toggle_10382_reset),
    .valid(toggle_10382_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(10446)) toggle_10446 (
    .clock(toggle_10446_clock),
    .reset(toggle_10446_reset),
    .valid(toggle_10446_valid)
  );
  GEN_w16_toggle #(.COVER_INDEX(10510)) toggle_10510 (
    .clock(toggle_10510_clock),
    .reset(toggle_10510_reset),
    .valid(toggle_10510_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10526)) toggle_10526 (
    .clock(toggle_10526_clock),
    .reset(toggle_10526_reset),
    .valid(toggle_10526_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10527)) toggle_10527 (
    .clock(toggle_10527_clock),
    .reset(toggle_10527_reset),
    .valid(toggle_10527_valid)
  );
  assign io__in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io__in_w_ready = io__in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io__in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io__in_ar_ready = io__in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io__in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io__in_r_bits_data = _io_in_r_bits_data_T_12 | _io_in_r_bits_data_T_9; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io__extra_mtip = io_extra_mtip_REG; // @[src/main/scala/device/AXI4CLINT.scala 66:21]
  assign io__extra_msip = io_extra_msip_REG; // @[src/main/scala/device/AXI4CLINT.scala 67:21]
  assign io_extra_mtip = io__extra_mtip;
  assign io_extra_msip = io__extra_msip;
  assign toggle_10185_clock = clock;
  assign toggle_10185_reset = reset;
  assign toggle_10185_valid = r_busy ^ toggle_10185_valid_reg;
  assign toggle_10186_clock = clock;
  assign toggle_10186_reset = reset;
  assign toggle_10186_valid = ren_REG ^ toggle_10186_valid_reg;
  assign toggle_10187_clock = clock;
  assign toggle_10187_reset = reset;
  assign toggle_10187_valid = io_in_r_valid_r ^ toggle_10187_valid_reg;
  assign toggle_10188_clock = clock;
  assign toggle_10188_reset = reset;
  assign toggle_10188_valid = w_busy ^ toggle_10188_valid_reg;
  assign toggle_10189_clock = clock;
  assign toggle_10189_reset = reset;
  assign toggle_10189_valid = io_in_b_valid_r ^ toggle_10189_valid_reg;
  assign toggle_10190_clock = clock;
  assign toggle_10190_reset = reset;
  assign toggle_10190_valid = mtime ^ toggle_10190_valid_reg;
  assign toggle_10254_clock = clock;
  assign toggle_10254_reset = reset;
  assign toggle_10254_valid = mtimecmp ^ toggle_10254_valid_reg;
  assign toggle_10318_clock = clock;
  assign toggle_10318_reset = reset;
  assign toggle_10318_valid = msip ^ toggle_10318_valid_reg;
  assign toggle_10382_clock = clock;
  assign toggle_10382_reset = reset;
  assign toggle_10382_valid = freq_reg ^ toggle_10382_valid_reg;
  assign toggle_10446_clock = clock;
  assign toggle_10446_reset = reset;
  assign toggle_10446_valid = inc_reg ^ toggle_10446_valid_reg;
  assign toggle_10510_clock = clock;
  assign toggle_10510_reset = reset;
  assign toggle_10510_valid = cnt ^ toggle_10510_valid_reg;
  assign toggle_10526_clock = clock;
  assign toggle_10526_reset = reset;
  assign toggle_10526_valid = io_extra_mtip_REG ^ toggle_10526_valid_reg;
  assign toggle_10527_clock = clock;
  assign toggle_10527_reset = reset;
  assign toggle_10527_valid = io_extra_msip_REG ^ toggle_10527_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 32:22]
      mtime <= 64'h0; // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'hbff8) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      mtime <= _mtime_T_7; // @[src/main/scala/utils/RegMap.scala 32:52]
    end else if (isWFI_0) begin // @[src/main/scala/device/AXI4CLINT.scala 51:18]
      mtime <= _mtime_T_3; // @[src/main/scala/device/AXI4CLINT.scala 51:26]
    end else if (tick) begin // @[src/main/scala/device/AXI4CLINT.scala 46:15]
      mtime <= _mtime_T_1; // @[src/main/scala/device/AXI4CLINT.scala 46:23]
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 33:25]
      mtimecmp <= 64'h0; // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'h4000) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      mtimecmp <= _mtimecmp_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 34:21]
      msip <= 64'h0; // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      msip <= _msip_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 37:25]
      freq_reg <= 64'h2710; // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'h8000) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      freq_reg <= _freq_reg_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 39:24]
      inc_reg <= 64'h1; // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[15:0] == 16'h8008) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      inc_reg <= _inc_reg_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4CLINT.scala 42:20]
      cnt <= 16'h0; // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    end else if (nextCnt < freq) begin // @[src/main/scala/device/AXI4CLINT.scala 44:13]
      cnt <= nextCnt;
    end else begin
      cnt <= 16'h0;
    end
    io_extra_mtip_REG <= mtime >= mtimecmp; // @[src/main/scala/device/AXI4CLINT.scala 66:38]
    io_extra_msip_REG <= msip != 64'h0; // @[src/main/scala/device/AXI4CLINT.scala 67:37]
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    r_busy_p <= r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10185_valid_reg <= r_busy;
    ren_REG_p <= ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    toggle_10186_valid_reg <= ren_REG;
    io_in_r_valid_r_p <= io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10187_valid_reg <= io_in_r_valid_r;
    w_busy_p <= w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10188_valid_reg <= w_busy;
    io_in_b_valid_r_p <= io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10189_valid_reg <= io_in_b_valid_r;
    mtime_p <= mtime; // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    toggle_10190_valid_reg <= mtime;
    mtimecmp_p <= mtimecmp; // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    toggle_10254_valid_reg <= mtimecmp;
    msip_p <= msip; // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    toggle_10318_valid_reg <= msip;
    freq_reg_p <= freq_reg; // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    toggle_10382_valid_reg <= freq_reg;
    inc_reg_p <= inc_reg; // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    toggle_10446_valid_reg <= inc_reg;
    cnt_p <= cnt; // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    toggle_10510_valid_reg <= cnt;
    io_extra_mtip_REG_p <= io_extra_mtip_REG; // @[src/main/scala/device/AXI4CLINT.scala 66:31]
    toggle_10526_valid_reg <= io_extra_mtip_REG;
    io_extra_msip_REG_p <= io_extra_msip_REG; // @[src/main/scala/device/AXI4CLINT.scala 67:31]
    toggle_10527_valid_reg <= io_extra_msip_REG;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  mtime = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mtimecmp = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  msip = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  freq_reg = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  inc_reg = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  cnt = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  io_extra_mtip_REG = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  io_extra_msip_REG = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  r_busy_p = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  toggle_10185_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  ren_REG_p = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  toggle_10186_valid_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  io_in_r_valid_r_p = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  toggle_10187_valid_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  w_busy_p = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  toggle_10188_valid_reg = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  io_in_b_valid_r_p = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  toggle_10189_valid_reg = _RAND_22[0:0];
  _RAND_23 = {2{`RANDOM}};
  mtime_p = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  toggle_10190_valid_reg = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  mtimecmp_p = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  toggle_10254_valid_reg = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  msip_p = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  toggle_10318_valid_reg = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  freq_reg_p = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  toggle_10382_valid_reg = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  inc_reg_p = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  toggle_10446_valid_reg = _RAND_32[63:0];
  _RAND_33 = {1{`RANDOM}};
  cnt_p = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  toggle_10510_valid_reg = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  io_extra_mtip_REG_p = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  toggle_10526_valid_reg = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  io_extra_msip_REG_p = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  toggle_10527_valid_reg = _RAND_38[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(r_busy_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(ren_REG_t); // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_valid_r_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(w_busy_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(io_in_b_valid_r_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[0]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[1]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[2]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[3]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[4]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[5]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[6]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[7]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[8]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[9]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[10]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[11]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[12]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[13]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[14]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[15]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[16]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[17]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[18]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[19]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[20]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[21]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[22]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[23]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[24]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[25]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[26]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[27]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[28]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[29]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[30]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[31]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[32]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[33]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[34]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[35]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[36]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[37]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[38]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[39]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[40]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[41]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[42]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[43]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[44]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[45]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[46]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[47]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[48]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[49]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[50]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[51]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[52]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[53]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[54]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[55]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[56]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[57]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[58]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[59]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[60]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[61]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[62]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtime_t[63]); // @[src/main/scala/device/AXI4CLINT.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[0]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[1]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[2]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[3]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[4]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[5]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[6]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[7]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[8]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[9]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[10]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[11]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[12]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[13]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[14]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[15]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[16]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[17]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[18]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[19]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[20]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[21]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[22]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[23]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[24]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[25]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[26]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[27]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[28]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[29]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[30]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[31]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[32]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[33]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[34]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[35]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[36]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[37]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[38]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[39]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[40]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[41]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[42]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[43]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[44]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[45]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[46]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[47]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[48]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[49]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[50]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[51]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[52]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[53]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[54]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[55]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[56]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[57]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[58]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[59]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[60]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[61]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[62]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(mtimecmp_t[63]); // @[src/main/scala/device/AXI4CLINT.scala 33:25]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[0]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[1]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[2]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[3]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[4]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[5]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[6]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[7]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[8]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[9]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[10]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[11]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[12]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[13]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[14]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[15]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[16]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[17]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[18]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[19]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[20]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[21]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[22]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[23]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[24]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[25]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[26]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[27]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[28]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[29]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[30]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[31]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[32]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[33]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[34]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[35]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[36]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[37]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[38]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[39]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[40]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[41]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[42]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[43]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[44]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[45]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[46]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[47]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[48]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[49]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[50]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[51]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[52]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[53]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[54]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[55]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[56]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[57]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[58]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[59]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[60]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[61]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[62]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(msip_t[63]); // @[src/main/scala/device/AXI4CLINT.scala 34:21]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[0]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[1]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[2]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[3]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[4]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[5]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[6]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[7]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[8]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[9]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[10]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[11]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[12]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[13]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[14]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[15]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[16]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[17]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[18]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[19]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[20]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[21]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[22]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[23]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[24]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[25]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[26]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[27]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[28]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[29]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[30]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[31]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[32]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[33]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[34]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[35]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[36]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[37]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[38]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[39]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[40]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[41]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[42]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[43]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[44]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[45]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[46]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[47]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[48]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[49]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[50]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[51]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[52]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[53]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[54]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[55]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[56]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[57]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[58]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[59]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[60]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[61]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[62]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(freq_reg_t[63]); // @[src/main/scala/device/AXI4CLINT.scala 37:25]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[0]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[1]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[2]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[3]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[4]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[5]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[6]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[7]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[8]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[9]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[10]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[11]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[12]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[13]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[14]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[15]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[16]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[17]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[18]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[19]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[20]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[21]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[22]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[23]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[24]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[25]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[26]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[27]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[28]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[29]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[30]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[31]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[32]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[33]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[34]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[35]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[36]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[37]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[38]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[39]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[40]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[41]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[42]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[43]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[44]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[45]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[46]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[47]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[48]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[49]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[50]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[51]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[52]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[53]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[54]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[55]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[56]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[57]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[58]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[59]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[60]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[61]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[62]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(inc_reg_t[63]); // @[src/main/scala/device/AXI4CLINT.scala 39:24]
    end
    //
    if (enToggle_past) begin
      cover(cnt_t[0]); // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    end
    //
    if (enToggle_past) begin
      cover(cnt_t[1]); // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    end
    //
    if (enToggle_past) begin
      cover(cnt_t[2]); // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    end
    //
    if (enToggle_past) begin
      cover(cnt_t[3]); // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    end
    //
    if (enToggle_past) begin
      cover(cnt_t[4]); // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    end
    //
    if (enToggle_past) begin
      cover(cnt_t[5]); // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    end
    //
    if (enToggle_past) begin
      cover(cnt_t[6]); // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    end
    //
    if (enToggle_past) begin
      cover(cnt_t[7]); // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    end
    //
    if (enToggle_past) begin
      cover(cnt_t[8]); // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    end
    //
    if (enToggle_past) begin
      cover(cnt_t[9]); // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    end
    //
    if (enToggle_past) begin
      cover(cnt_t[10]); // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    end
    //
    if (enToggle_past) begin
      cover(cnt_t[11]); // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    end
    //
    if (enToggle_past) begin
      cover(cnt_t[12]); // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    end
    //
    if (enToggle_past) begin
      cover(cnt_t[13]); // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    end
    //
    if (enToggle_past) begin
      cover(cnt_t[14]); // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    end
    //
    if (enToggle_past) begin
      cover(cnt_t[15]); // @[src/main/scala/device/AXI4CLINT.scala 42:20]
    end
    //
    if (enToggle_past) begin
      cover(io_extra_mtip_REG_t); // @[src/main/scala/device/AXI4CLINT.scala 66:31]
    end
    //
    if (enToggle_past) begin
      cover(io_extra_msip_REG_t); // @[src/main/scala/device/AXI4CLINT.scala 67:31]
    end
  end
endmodule
module SimpleBus2AXI4Converter_1(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_resp_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_aw_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_out_w_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_w_bits_strb, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_b_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_ar_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_r_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_out_r_bits_data // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  toAXI4Lite = ~(io_in_req_valid & io_in_req_bits_cmd[1]); // @[src/main/scala/bus/simplebus/ToAXI4.scala 151:20]
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 | awAck & wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 189:53]
  wire  _GEN_2 = _wSend_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wen_T_1 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  _io_out_ar_valid_T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _io_out_aw_valid_T_1 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  wire  _io_out_w_valid_T_2 = ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:36]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  awAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  awAck_t = awAck ^ awAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10528_clock;
  wire  toggle_10528_reset;
  wire  toggle_10528_valid;
  reg  toggle_10528_valid_reg;
  reg  wAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wAck_t = wAck ^ wAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10529_clock;
  wire  toggle_10529_reset;
  wire  toggle_10529_valid;
  reg  toggle_10529_valid_reg;
  reg  wen_p; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  wen_t = wen ^ wen_p; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  toggle_10530_clock;
  wire  toggle_10530_reset;
  wire  toggle_10530_valid;
  reg  toggle_10530_valid_reg;
  GEN_w1_toggle #(.COVER_INDEX(10528)) toggle_10528 (
    .clock(toggle_10528_clock),
    .reset(toggle_10528_reset),
    .valid(toggle_10528_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10529)) toggle_10529 (
    .clock(toggle_10529_clock),
    .reset(toggle_10529_reset),
    .valid(toggle_10529_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10530)) toggle_10530 (
    .clock(toggle_10530_clock),
    .reset(toggle_10530_reset),
    .valid(toggle_10530_valid)
  );
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _io_out_w_valid_T_2 & io_out_w_ready : io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 199:25]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 183:23]
  assign io_out_aw_valid = _io_out_aw_valid_T_1 & ~awAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 193:33]
  assign io_out_aw_bits_addr = io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_w_valid = _io_out_aw_valid_T_1 & ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:33]
  assign io_out_w_bits_data = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 160:10]
  assign io_out_w_bits_strb = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 161:10]
  assign io_out_b_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 198:16]
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 158:12]
  assign io_out_r_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 197:16]
  assign toggle_10528_clock = clock;
  assign toggle_10528_reset = reset;
  assign toggle_10528_valid = awAck ^ toggle_10528_valid_reg;
  assign toggle_10529_clock = clock;
  assign toggle_10529_reset = reset;
  assign toggle_10529_valid = wAck ^ toggle_10529_valid_reg;
  assign toggle_10530_clock = clock;
  assign toggle_10530_reset = reset;
  assign toggle_10530_valid = wen ^ toggle_10530_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_2;
    end
    if (_wen_T_1) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
      wen <= io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~toAXI4Lite) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    awAck_p <= awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10528_valid_reg <= awAck;
    wAck_p <= wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10529_valid_reg <= wAck;
    wen_p <= wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    toggle_10530_valid_reg <= wen;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  awAck_p = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  toggle_10528_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  wAck_p = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  toggle_10529_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  wen_p = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  toggle_10530_valid_reg = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(toAXI4Lite); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
    end
    //
    if (enToggle_past) begin
      cover(awAck_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(wAck_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(wen_t); // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
  end
endmodule
module AXI4PLIC(
  input         clock,
  input         reset,
  output        io__in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io__in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io__in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io__in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io__in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io__in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io__in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io__extra_meip_0, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_meip_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  wire  _r_busy_T = io__in_ar_ready & io__in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _r_busy_T_1 = io__in_r_ready & io__in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _r_busy_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_2 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io__in_aw_ready & io__in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io__in_b_ready & io__in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _w_busy_T | _GEN_4; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io__in_w_ready & io__in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [31:0] priority_0; // @[src/main/scala/device/AXI4PLIC.scala 37:39]
  reg [31:0] enable_0_0; // @[src/main/scala/device/AXI4PLIC.scala 48:64]
  reg [31:0] threshold_0; // @[src/main/scala/device/AXI4PLIC.scala 53:40]
  wire [7:0] _T_12 = io__in_w_bits_strb >> io__in_aw_bits_addr[2:0]; // @[src/main/scala/device/AXI4PLIC.scala 89:85]
  wire [7:0] _T_21 = _T_12[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_22 = _T_12[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_23 = _T_12[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_24 = _T_12[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_25 = _T_12[4] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_26 = _T_12[5] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_27 = _T_12[6] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_28 = _T_12[7] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [63:0] _T_29 = {_T_28,_T_27,_T_26,_T_25,_T_24,_T_23,_T_22,_T_21}; // @[src/main/scala/utils/BitUtils.scala 27:27]
  wire  _rdata_T_1 = 26'h2000 == io__in_ar_bits_addr[25:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_3 = 26'h4 == io__in_ar_bits_addr[25:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_4 = 26'h200000 == io__in_ar_bits_addr[25:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _rdata_T_6 = _rdata_T_1 ? enable_0_0 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_8 = _rdata_T_3 ? priority_0 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_9 = _rdata_T_4 ? threshold_0 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_12 = _rdata_T_6 | _rdata_T_8; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] rdata = _rdata_T_12 | _rdata_T_9; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _enable_0_0_T = io__in_w_bits_data[31:0] & _T_29[31:0]; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [31:0] _enable_0_0_T_1 = ~_T_29[31:0]; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [31:0] _enable_0_0_T_2 = enable_0_0 & _enable_0_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _enable_0_0_T_3 = _enable_0_0_T | _enable_0_0_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _priority_0_T_2 = priority_0 & _enable_0_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _priority_0_T_3 = _enable_0_0_T | _priority_0_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _threshold_0_T_2 = threshold_0 & _enable_0_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _threshold_0_T_3 = _enable_0_0_T | _threshold_0_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  r_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  r_busy_t = r_busy ^ r_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10531_clock;
  wire  toggle_10531_reset;
  wire  toggle_10531_valid;
  reg  toggle_10531_valid_reg;
  reg  ren_REG_p; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  ren_REG_t = ren_REG ^ ren_REG_p; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  toggle_10532_clock;
  wire  toggle_10532_reset;
  wire  toggle_10532_valid;
  reg  toggle_10532_valid_reg;
  reg  io_in_r_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  io_in_r_valid_r_t = io_in_r_valid_r ^ io_in_r_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10533_clock;
  wire  toggle_10533_reset;
  wire  toggle_10533_valid;
  reg  toggle_10533_valid_reg;
  reg  w_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  w_busy_t = w_busy ^ w_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10534_clock;
  wire  toggle_10534_reset;
  wire  toggle_10534_valid;
  reg  toggle_10534_valid_reg;
  reg  io_in_b_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  io_in_b_valid_r_t = io_in_b_valid_r ^ io_in_b_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10535_clock;
  wire  toggle_10535_reset;
  wire  toggle_10535_valid;
  reg  toggle_10535_valid_reg;
  reg [31:0] priority_0_p; // @[src/main/scala/device/AXI4PLIC.scala 37:39]
  wire [31:0] priority_0_t = priority_0 ^ priority_0_p; // @[src/main/scala/device/AXI4PLIC.scala 37:39]
  wire  toggle_10536_clock;
  wire  toggle_10536_reset;
  wire [31:0] toggle_10536_valid;
  reg [31:0] toggle_10536_valid_reg;
  reg [31:0] enable_0_0_p; // @[src/main/scala/device/AXI4PLIC.scala 48:64]
  wire [31:0] enable_0_0_t = enable_0_0 ^ enable_0_0_p; // @[src/main/scala/device/AXI4PLIC.scala 48:64]
  wire  toggle_10568_clock;
  wire  toggle_10568_reset;
  wire [31:0] toggle_10568_valid;
  reg [31:0] toggle_10568_valid_reg;
  reg [31:0] threshold_0_p; // @[src/main/scala/device/AXI4PLIC.scala 53:40]
  wire [31:0] threshold_0_t = threshold_0 ^ threshold_0_p; // @[src/main/scala/device/AXI4PLIC.scala 53:40]
  wire  toggle_10600_clock;
  wire  toggle_10600_reset;
  wire [31:0] toggle_10600_valid;
  reg [31:0] toggle_10600_valid_reg;
  GEN_w1_toggle #(.COVER_INDEX(10531)) toggle_10531 (
    .clock(toggle_10531_clock),
    .reset(toggle_10531_reset),
    .valid(toggle_10531_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10532)) toggle_10532 (
    .clock(toggle_10532_clock),
    .reset(toggle_10532_reset),
    .valid(toggle_10532_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10533)) toggle_10533 (
    .clock(toggle_10533_clock),
    .reset(toggle_10533_reset),
    .valid(toggle_10533_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10534)) toggle_10534 (
    .clock(toggle_10534_clock),
    .reset(toggle_10534_reset),
    .valid(toggle_10534_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10535)) toggle_10535 (
    .clock(toggle_10535_clock),
    .reset(toggle_10535_reset),
    .valid(toggle_10535_valid)
  );
  GEN_w32_toggle #(.COVER_INDEX(10536)) toggle_10536 (
    .clock(toggle_10536_clock),
    .reset(toggle_10536_reset),
    .valid(toggle_10536_valid)
  );
  GEN_w32_toggle #(.COVER_INDEX(10568)) toggle_10568 (
    .clock(toggle_10568_clock),
    .reset(toggle_10568_reset),
    .valid(toggle_10568_valid)
  );
  GEN_w32_toggle #(.COVER_INDEX(10600)) toggle_10600 (
    .clock(toggle_10600_clock),
    .reset(toggle_10600_reset),
    .valid(toggle_10600_valid)
  );
  assign io__in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io__in_w_ready = io__in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io__in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io__in_ar_ready = io__in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io__in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io__in_r_bits_data = {rdata,rdata}; // @[src/main/scala/device/AXI4PLIC.scala 91:25]
  assign io__extra_meip_0 = 1'h0; // @[src/main/scala/device/AXI4PLIC.scala 93:87]
  assign io_extra_meip_0 = io__extra_meip_0;
  assign toggle_10531_clock = clock;
  assign toggle_10531_reset = reset;
  assign toggle_10531_valid = r_busy ^ toggle_10531_valid_reg;
  assign toggle_10532_clock = clock;
  assign toggle_10532_reset = reset;
  assign toggle_10532_valid = ren_REG ^ toggle_10532_valid_reg;
  assign toggle_10533_clock = clock;
  assign toggle_10533_reset = reset;
  assign toggle_10533_valid = io_in_r_valid_r ^ toggle_10533_valid_reg;
  assign toggle_10534_clock = clock;
  assign toggle_10534_reset = reset;
  assign toggle_10534_valid = w_busy ^ toggle_10534_valid_reg;
  assign toggle_10535_clock = clock;
  assign toggle_10535_reset = reset;
  assign toggle_10535_valid = io_in_b_valid_r ^ toggle_10535_valid_reg;
  assign toggle_10536_clock = clock;
  assign toggle_10536_reset = reset;
  assign toggle_10536_valid = priority_0 ^ toggle_10536_valid_reg;
  assign toggle_10568_clock = clock;
  assign toggle_10568_reset = reset;
  assign toggle_10568_valid = enable_0_0 ^ toggle_10568_valid_reg;
  assign toggle_10600_clock = clock;
  assign toggle_10600_reset = reset;
  assign toggle_10600_valid = threshold_0 ^ toggle_10600_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
    if (_io_in_b_valid_T & io__in_aw_bits_addr[25:0] == 26'h4) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      priority_0 <= _priority_0_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4PLIC.scala 48:64]
      enable_0_0 <= 32'h0; // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end else if (_io_in_b_valid_T & io__in_aw_bits_addr[25:0] == 26'h2000) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      enable_0_0 <= _enable_0_0_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (_io_in_b_valid_T & io__in_aw_bits_addr[25:0] == 26'h200000) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      threshold_0 <= _threshold_0_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    r_busy_p <= r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10531_valid_reg <= r_busy;
    ren_REG_p <= ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    toggle_10532_valid_reg <= ren_REG;
    io_in_r_valid_r_p <= io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10533_valid_reg <= io_in_r_valid_r;
    w_busy_p <= w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10534_valid_reg <= w_busy;
    io_in_b_valid_r_p <= io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10535_valid_reg <= io_in_b_valid_r;
    priority_0_p <= priority_0; // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    toggle_10536_valid_reg <= priority_0;
    enable_0_0_p <= enable_0_0; // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    toggle_10568_valid_reg <= enable_0_0;
    threshold_0_p <= threshold_0; // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    toggle_10600_valid_reg <= threshold_0;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  priority_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  enable_0_0 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  threshold_0 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  r_busy_p = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  toggle_10531_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ren_REG_p = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  toggle_10532_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  io_in_r_valid_r_p = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  toggle_10533_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  w_busy_p = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  toggle_10534_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  io_in_b_valid_r_p = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  toggle_10535_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  priority_0_p = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  toggle_10536_valid_reg = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  enable_0_0_p = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  toggle_10568_valid_reg = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  threshold_0_p = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  toggle_10600_valid_reg = _RAND_23[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(r_busy_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(ren_REG_t); // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_valid_r_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(w_busy_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(io_in_b_valid_r_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[0]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[1]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[2]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[3]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[4]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[5]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[6]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[7]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[8]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[9]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[10]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[11]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[12]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[13]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[14]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[15]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[16]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[17]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[18]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[19]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[20]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[21]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[22]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[23]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[24]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[25]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[26]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[27]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[28]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[29]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[30]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(priority_0_t[31]); // @[src/main/scala/device/AXI4PLIC.scala 37:39]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[0]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[1]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[2]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[3]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[4]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[5]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[6]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[7]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[8]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[9]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[10]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[11]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[12]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[13]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[14]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[15]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[16]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[17]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[18]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[19]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[20]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[21]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[22]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[23]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[24]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[25]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[26]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[27]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[28]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[29]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[30]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(enable_0_0_t[31]); // @[src/main/scala/device/AXI4PLIC.scala 48:64]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[0]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[1]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[2]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[3]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[4]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[5]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[6]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[7]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[8]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[9]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[10]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[11]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[12]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[13]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[14]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[15]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[16]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[17]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[18]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[19]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[20]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[21]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[22]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[23]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[24]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[25]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[26]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[27]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[28]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[29]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[30]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
    //
    if (enToggle_past) begin
      cover(threshold_0_t[31]); // @[src/main/scala/device/AXI4PLIC.scala 53:40]
    end
  end
endmodule
module SimpleBus2AXI4Converter_2(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_resp_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_aw_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_out_w_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_w_bits_strb, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_b_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_ar_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_r_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_out_r_bits_data // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  toAXI4Lite = ~(io_in_req_valid & io_in_req_bits_cmd[1]); // @[src/main/scala/bus/simplebus/ToAXI4.scala 151:20]
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 | awAck & wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 189:53]
  wire  _GEN_2 = _wSend_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wen_T_1 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  _io_out_ar_valid_T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _io_out_aw_valid_T_1 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  wire  _io_out_w_valid_T_2 = ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:36]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  awAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  awAck_t = awAck ^ awAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10632_clock;
  wire  toggle_10632_reset;
  wire  toggle_10632_valid;
  reg  toggle_10632_valid_reg;
  reg  wAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wAck_t = wAck ^ wAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10633_clock;
  wire  toggle_10633_reset;
  wire  toggle_10633_valid;
  reg  toggle_10633_valid_reg;
  reg  wen_p; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  wen_t = wen ^ wen_p; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  toggle_10634_clock;
  wire  toggle_10634_reset;
  wire  toggle_10634_valid;
  reg  toggle_10634_valid_reg;
  GEN_w1_toggle #(.COVER_INDEX(10632)) toggle_10632 (
    .clock(toggle_10632_clock),
    .reset(toggle_10632_reset),
    .valid(toggle_10632_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10633)) toggle_10633 (
    .clock(toggle_10633_clock),
    .reset(toggle_10633_reset),
    .valid(toggle_10633_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10634)) toggle_10634 (
    .clock(toggle_10634_clock),
    .reset(toggle_10634_reset),
    .valid(toggle_10634_valid)
  );
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _io_out_w_valid_T_2 & io_out_w_ready : io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 199:25]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 183:23]
  assign io_out_aw_valid = _io_out_aw_valid_T_1 & ~awAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 193:33]
  assign io_out_aw_bits_addr = io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_w_valid = _io_out_aw_valid_T_1 & ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:33]
  assign io_out_w_bits_data = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 160:10]
  assign io_out_w_bits_strb = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 161:10]
  assign io_out_b_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 198:16]
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 158:12]
  assign io_out_r_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 197:16]
  assign toggle_10632_clock = clock;
  assign toggle_10632_reset = reset;
  assign toggle_10632_valid = awAck ^ toggle_10632_valid_reg;
  assign toggle_10633_clock = clock;
  assign toggle_10633_reset = reset;
  assign toggle_10633_valid = wAck ^ toggle_10633_valid_reg;
  assign toggle_10634_clock = clock;
  assign toggle_10634_reset = reset;
  assign toggle_10634_valid = wen ^ toggle_10634_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_2;
    end
    if (_wen_T_1) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
      wen <= io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~toAXI4Lite) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    awAck_p <= awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10632_valid_reg <= awAck;
    wAck_p <= wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10633_valid_reg <= wAck;
    wen_p <= wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    toggle_10634_valid_reg <= wen;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  awAck_p = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  toggle_10632_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  wAck_p = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  toggle_10633_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  wen_p = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  toggle_10634_valid_reg = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(toAXI4Lite); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
    end
    //
    if (enToggle_past) begin
      cover(awAck_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(wAck_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(wen_t); // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
  end
endmodule
module NutShell(
  input         clock,
  input         reset,
  input         io_mem_aw_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mem_aw_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  output [31:0] io_mem_aw_bits_addr, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mem_w_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mem_w_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  output [63:0] io_mem_w_bits_data, // @[src/main/scala/system/NutShell.scala 45:14]
  output [7:0]  io_mem_w_bits_strb, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mem_w_bits_last, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mem_b_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mem_ar_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  output [31:0] io_mem_ar_bits_addr, // @[src/main/scala/system/NutShell.scala 45:14]
  output [7:0]  io_mem_ar_bits_len, // @[src/main/scala/system/NutShell.scala 45:14]
  output [2:0]  io_mem_ar_bits_size, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mem_r_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  input  [63:0] io_mem_r_bits_data, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mem_r_bits_last, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mmio_req_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mmio_req_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  output [31:0] io_mmio_req_bits_addr, // @[src/main/scala/system/NutShell.scala 45:14]
  output [3:0]  io_mmio_req_bits_cmd, // @[src/main/scala/system/NutShell.scala 45:14]
  output [7:0]  io_mmio_req_bits_wmask, // @[src/main/scala/system/NutShell.scala 45:14]
  output [63:0] io_mmio_req_bits_wdata, // @[src/main/scala/system/NutShell.scala 45:14]
  output        io_mmio_resp_ready, // @[src/main/scala/system/NutShell.scala 45:14]
  input         io_mmio_resp_valid, // @[src/main/scala/system/NutShell.scala 45:14]
  input  [3:0]  io_mmio_resp_bits_cmd, // @[src/main/scala/system/NutShell.scala 45:14]
  input  [63:0] io_mmio_resp_bits_rdata // @[src/main/scala/system/NutShell.scala 45:14]
);
  wire  nutcore_clock; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_reset; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_req_ready; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_req_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [31:0] nutcore_io_imem_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_resp_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_imem_mem_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_req_ready; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_req_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [31:0] nutcore_io_dmem_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [2:0] nutcore_io_dmem_mem_req_bits_size; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_mem_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [7:0] nutcore_io_dmem_mem_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_mem_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_resp_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_mem_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_mem_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_mmio_req_ready; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_mmio_req_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [31:0] nutcore_io_mmio_req_bits_addr; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_mmio_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [7:0] nutcore_io_mmio_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_mmio_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_mmio_resp_valid; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [3:0] nutcore_io_mmio_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 53:23]
  wire [63:0] nutcore_io_mmio_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_extra_meip_0; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_isWFI; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_extra_mtip; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  nutcore_io_extra_msip; // @[src/main/scala/system/NutShell.scala 53:23]
  wire  cohMg_clock; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_reset; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_in_req_valid; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [31:0] cohMg_io_in_req_bits_addr; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [3:0] cohMg_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [63:0] cohMg_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_out_mem_req_ready; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_out_mem_req_valid; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [31:0] cohMg_io_out_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_out_mem_resp_ready; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  cohMg_io_out_mem_resp_valid; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [3:0] cohMg_io_out_mem_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_mem_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 54:21]
  wire  xbar_clock; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_reset; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_0_req_ready; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_0_req_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [31:0] xbar_io_in_0_req_bits_addr; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_0_resp_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_in_0_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_in_0_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_1_req_ready; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_1_req_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [31:0] xbar_io_in_1_req_bits_addr; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [2:0] xbar_io_in_1_req_bits_size; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_in_1_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [7:0] xbar_io_in_1_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_in_1_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_in_1_resp_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_in_1_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_in_1_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_out_req_ready; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_out_req_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [31:0] xbar_io_out_req_bits_addr; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [2:0] xbar_io_out_req_bits_size; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_out_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [7:0] xbar_io_out_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_out_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_out_resp_ready; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  xbar_io_out_resp_valid; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [3:0] xbar_io_out_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 55:20]
  wire [63:0] xbar_io_out_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 55:20]
  wire  axi2sb_clock; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  axi2sb_reset; // @[src/main/scala/system/NutShell.scala 61:22]
  wire  memport_bridge_clock; // @[src/main/scala/bus/simplebus/ToMemPort.scala 50:24]
  wire  memport_bridge_reset; // @[src/main/scala/bus/simplebus/ToMemPort.scala 50:24]
  wire  memAddrMap_clock; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_reset; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_in_req_valid; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [31:0] memAddrMap_io_in_req_bits_addr; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [2:0] memAddrMap_io_in_req_bits_size; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_in_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [7:0] memAddrMap_io_in_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_in_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_out_req_ready; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_out_req_valid; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [31:0] memAddrMap_io_out_req_bits_addr; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [2:0] memAddrMap_io_out_req_bits_size; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_out_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [7:0] memAddrMap_io_out_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_out_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  memAddrMap_io_out_resp_valid; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_out_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_out_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 93:26]
  wire  io_mem_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] io_mem_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [2:0] io_mem_bridge_io_in_req_bits_size; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] io_mem_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] io_mem_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] io_mem_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] io_mem_bridge_io_in_resp_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] io_mem_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] io_mem_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] io_mem_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] io_mem_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_w_bits_last; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] io_mem_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] io_mem_bridge_io_out_ar_bits_len; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [2:0] io_mem_bridge_io_out_ar_bits_size; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] io_mem_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  io_mem_bridge_io_out_r_bits_last; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  mmioXbar_clock; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_reset; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_in_req_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_in_req_bits_addr; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_in_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_in_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_in_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_req_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_req_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_0_req_bits_addr; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_0_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_0_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_0_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_resp_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_resp_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_0_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_req_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_req_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_1_req_bits_addr; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_1_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_1_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_1_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_resp_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_resp_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_1_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_req_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_req_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_2_req_bits_addr; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_2_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_2_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_2_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_resp_ready; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_resp_valid; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_2_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_2_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 106:24]
  wire  clint_clock; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_reset; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_aw_ready; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_aw_valid; // @[src/main/scala/system/NutShell.scala 113:21]
  wire [31:0] clint_io__in_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_w_ready; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_w_valid; // @[src/main/scala/system/NutShell.scala 113:21]
  wire [63:0] clint_io__in_w_bits_data; // @[src/main/scala/system/NutShell.scala 113:21]
  wire [7:0] clint_io__in_w_bits_strb; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_b_ready; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_b_valid; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_ar_ready; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_ar_valid; // @[src/main/scala/system/NutShell.scala 113:21]
  wire [31:0] clint_io__in_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_r_ready; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__in_r_valid; // @[src/main/scala/system/NutShell.scala 113:21]
  wire [63:0] clint_io__in_r_bits_data; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__extra_mtip; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io__extra_msip; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_isWFI_0; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io_extra_mtip; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io_extra_msip; // @[src/main/scala/system/NutShell.scala 113:21]
  wire  clint_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] clint_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] clint_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] clint_io_in_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] clint_io_in_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] clint_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] clint_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] clint_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] clint_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] clint_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  clint_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] clint_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_clock; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_reset; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_aw_ready; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_aw_valid; // @[src/main/scala/system/NutShell.scala 120:20]
  wire [31:0] plic_io__in_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_w_ready; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_w_valid; // @[src/main/scala/system/NutShell.scala 120:20]
  wire [63:0] plic_io__in_w_bits_data; // @[src/main/scala/system/NutShell.scala 120:20]
  wire [7:0] plic_io__in_w_bits_strb; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_b_ready; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_b_valid; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_ar_ready; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_ar_valid; // @[src/main/scala/system/NutShell.scala 120:20]
  wire [31:0] plic_io__in_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_r_ready; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__in_r_valid; // @[src/main/scala/system/NutShell.scala 120:20]
  wire [63:0] plic_io__in_r_bits_data; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io__extra_meip_0; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io_extra_meip_0; // @[src/main/scala/system/NutShell.scala 120:20]
  wire  plic_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] plic_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] plic_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] plic_io_in_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] plic_io_in_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] plic_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] plic_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] plic_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] plic_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] plic_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  plic_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] plic_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  NutCore nutcore ( // @[src/main/scala/system/NutShell.scala 53:23]
    .clock(nutcore_clock),
    .reset(nutcore_reset),
    .io_imem_mem_req_ready(nutcore_io_imem_mem_req_ready),
    .io_imem_mem_req_valid(nutcore_io_imem_mem_req_valid),
    .io_imem_mem_req_bits_addr(nutcore_io_imem_mem_req_bits_addr),
    .io_imem_mem_resp_valid(nutcore_io_imem_mem_resp_valid),
    .io_imem_mem_resp_bits_rdata(nutcore_io_imem_mem_resp_bits_rdata),
    .io_dmem_mem_req_ready(nutcore_io_dmem_mem_req_ready),
    .io_dmem_mem_req_valid(nutcore_io_dmem_mem_req_valid),
    .io_dmem_mem_req_bits_addr(nutcore_io_dmem_mem_req_bits_addr),
    .io_dmem_mem_req_bits_size(nutcore_io_dmem_mem_req_bits_size),
    .io_dmem_mem_req_bits_cmd(nutcore_io_dmem_mem_req_bits_cmd),
    .io_dmem_mem_req_bits_wmask(nutcore_io_dmem_mem_req_bits_wmask),
    .io_dmem_mem_req_bits_wdata(nutcore_io_dmem_mem_req_bits_wdata),
    .io_dmem_mem_resp_valid(nutcore_io_dmem_mem_resp_valid),
    .io_dmem_mem_resp_bits_cmd(nutcore_io_dmem_mem_resp_bits_cmd),
    .io_dmem_mem_resp_bits_rdata(nutcore_io_dmem_mem_resp_bits_rdata),
    .io_mmio_req_ready(nutcore_io_mmio_req_ready),
    .io_mmio_req_valid(nutcore_io_mmio_req_valid),
    .io_mmio_req_bits_addr(nutcore_io_mmio_req_bits_addr),
    .io_mmio_req_bits_cmd(nutcore_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(nutcore_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(nutcore_io_mmio_req_bits_wdata),
    .io_mmio_resp_valid(nutcore_io_mmio_resp_valid),
    .io_mmio_resp_bits_cmd(nutcore_io_mmio_resp_bits_cmd),
    .io_mmio_resp_bits_rdata(nutcore_io_mmio_resp_bits_rdata),
    .io_extra_meip_0(nutcore_io_extra_meip_0),
    .isWFI(nutcore_isWFI),
    .io_extra_mtip(nutcore_io_extra_mtip),
    .io_extra_msip(nutcore_io_extra_msip)
  );
  CoherenceManager cohMg ( // @[src/main/scala/system/NutShell.scala 54:21]
    .clock(cohMg_clock),
    .reset(cohMg_reset),
    .io_in_req_ready(cohMg_io_in_req_ready),
    .io_in_req_valid(cohMg_io_in_req_valid),
    .io_in_req_bits_addr(cohMg_io_in_req_bits_addr),
    .io_in_resp_valid(cohMg_io_in_resp_valid),
    .io_in_resp_bits_cmd(cohMg_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(cohMg_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(cohMg_io_out_mem_req_ready),
    .io_out_mem_req_valid(cohMg_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(cohMg_io_out_mem_req_bits_addr),
    .io_out_mem_resp_ready(cohMg_io_out_mem_resp_ready),
    .io_out_mem_resp_valid(cohMg_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(cohMg_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(cohMg_io_out_mem_resp_bits_rdata)
  );
  SimpleBusCrossbarNto1_2 xbar ( // @[src/main/scala/system/NutShell.scala 55:20]
    .clock(xbar_clock),
    .reset(xbar_reset),
    .io_in_0_req_ready(xbar_io_in_0_req_ready),
    .io_in_0_req_valid(xbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(xbar_io_in_0_req_bits_addr),
    .io_in_0_resp_valid(xbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_cmd(xbar_io_in_0_resp_bits_cmd),
    .io_in_0_resp_bits_rdata(xbar_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(xbar_io_in_1_req_ready),
    .io_in_1_req_valid(xbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(xbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_size(xbar_io_in_1_req_bits_size),
    .io_in_1_req_bits_cmd(xbar_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(xbar_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(xbar_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(xbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(xbar_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(xbar_io_in_1_resp_bits_rdata),
    .io_out_req_ready(xbar_io_out_req_ready),
    .io_out_req_valid(xbar_io_out_req_valid),
    .io_out_req_bits_addr(xbar_io_out_req_bits_addr),
    .io_out_req_bits_size(xbar_io_out_req_bits_size),
    .io_out_req_bits_cmd(xbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(xbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(xbar_io_out_req_bits_wdata),
    .io_out_resp_ready(xbar_io_out_resp_ready),
    .io_out_resp_valid(xbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(xbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(xbar_io_out_resp_bits_rdata)
  );
  AXI42SimpleBusConverter axi2sb ( // @[src/main/scala/system/NutShell.scala 61:22]
    .clock(axi2sb_clock),
    .reset(axi2sb_reset)
  );
  SimpleBus2MemPortConverter memport_bridge ( // @[src/main/scala/bus/simplebus/ToMemPort.scala 50:24]
    .clock(memport_bridge_clock),
    .reset(memport_bridge_reset)
  );
  SimpleBusAddressMapper memAddrMap ( // @[src/main/scala/system/NutShell.scala 93:26]
    .clock(memAddrMap_clock),
    .reset(memAddrMap_reset),
    .io_in_req_ready(memAddrMap_io_in_req_ready),
    .io_in_req_valid(memAddrMap_io_in_req_valid),
    .io_in_req_bits_addr(memAddrMap_io_in_req_bits_addr),
    .io_in_req_bits_size(memAddrMap_io_in_req_bits_size),
    .io_in_req_bits_cmd(memAddrMap_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(memAddrMap_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(memAddrMap_io_in_req_bits_wdata),
    .io_in_resp_valid(memAddrMap_io_in_resp_valid),
    .io_in_resp_bits_cmd(memAddrMap_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(memAddrMap_io_in_resp_bits_rdata),
    .io_out_req_ready(memAddrMap_io_out_req_ready),
    .io_out_req_valid(memAddrMap_io_out_req_valid),
    .io_out_req_bits_addr(memAddrMap_io_out_req_bits_addr),
    .io_out_req_bits_size(memAddrMap_io_out_req_bits_size),
    .io_out_req_bits_cmd(memAddrMap_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(memAddrMap_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(memAddrMap_io_out_req_bits_wdata),
    .io_out_resp_valid(memAddrMap_io_out_resp_valid),
    .io_out_resp_bits_cmd(memAddrMap_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(memAddrMap_io_out_resp_bits_rdata)
  );
  SimpleBus2AXI4Converter io_mem_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(io_mem_bridge_clock),
    .reset(io_mem_bridge_reset),
    .io_in_req_ready(io_mem_bridge_io_in_req_ready),
    .io_in_req_valid(io_mem_bridge_io_in_req_valid),
    .io_in_req_bits_addr(io_mem_bridge_io_in_req_bits_addr),
    .io_in_req_bits_size(io_mem_bridge_io_in_req_bits_size),
    .io_in_req_bits_cmd(io_mem_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(io_mem_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(io_mem_bridge_io_in_req_bits_wdata),
    .io_in_resp_valid(io_mem_bridge_io_in_resp_valid),
    .io_in_resp_bits_cmd(io_mem_bridge_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(io_mem_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(io_mem_bridge_io_out_aw_ready),
    .io_out_aw_valid(io_mem_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(io_mem_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(io_mem_bridge_io_out_w_ready),
    .io_out_w_valid(io_mem_bridge_io_out_w_valid),
    .io_out_w_bits_data(io_mem_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(io_mem_bridge_io_out_w_bits_strb),
    .io_out_w_bits_last(io_mem_bridge_io_out_w_bits_last),
    .io_out_b_valid(io_mem_bridge_io_out_b_valid),
    .io_out_ar_valid(io_mem_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(io_mem_bridge_io_out_ar_bits_addr),
    .io_out_ar_bits_len(io_mem_bridge_io_out_ar_bits_len),
    .io_out_ar_bits_size(io_mem_bridge_io_out_ar_bits_size),
    .io_out_r_valid(io_mem_bridge_io_out_r_valid),
    .io_out_r_bits_data(io_mem_bridge_io_out_r_bits_data),
    .io_out_r_bits_last(io_mem_bridge_io_out_r_bits_last)
  );
  SimpleBusCrossbar1toN mmioXbar ( // @[src/main/scala/system/NutShell.scala 106:24]
    .clock(mmioXbar_clock),
    .reset(mmioXbar_reset),
    .io_in_req_ready(mmioXbar_io_in_req_ready),
    .io_in_req_valid(mmioXbar_io_in_req_valid),
    .io_in_req_bits_addr(mmioXbar_io_in_req_bits_addr),
    .io_in_req_bits_cmd(mmioXbar_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(mmioXbar_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(mmioXbar_io_in_req_bits_wdata),
    .io_in_resp_valid(mmioXbar_io_in_resp_valid),
    .io_in_resp_bits_cmd(mmioXbar_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(mmioXbar_io_in_resp_bits_rdata),
    .io_out_0_req_ready(mmioXbar_io_out_0_req_ready),
    .io_out_0_req_valid(mmioXbar_io_out_0_req_valid),
    .io_out_0_req_bits_addr(mmioXbar_io_out_0_req_bits_addr),
    .io_out_0_req_bits_cmd(mmioXbar_io_out_0_req_bits_cmd),
    .io_out_0_req_bits_wmask(mmioXbar_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wdata(mmioXbar_io_out_0_req_bits_wdata),
    .io_out_0_resp_ready(mmioXbar_io_out_0_resp_ready),
    .io_out_0_resp_valid(mmioXbar_io_out_0_resp_valid),
    .io_out_0_resp_bits_rdata(mmioXbar_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(mmioXbar_io_out_1_req_ready),
    .io_out_1_req_valid(mmioXbar_io_out_1_req_valid),
    .io_out_1_req_bits_addr(mmioXbar_io_out_1_req_bits_addr),
    .io_out_1_req_bits_cmd(mmioXbar_io_out_1_req_bits_cmd),
    .io_out_1_req_bits_wmask(mmioXbar_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wdata(mmioXbar_io_out_1_req_bits_wdata),
    .io_out_1_resp_ready(mmioXbar_io_out_1_resp_ready),
    .io_out_1_resp_valid(mmioXbar_io_out_1_resp_valid),
    .io_out_1_resp_bits_rdata(mmioXbar_io_out_1_resp_bits_rdata),
    .io_out_2_req_ready(mmioXbar_io_out_2_req_ready),
    .io_out_2_req_valid(mmioXbar_io_out_2_req_valid),
    .io_out_2_req_bits_addr(mmioXbar_io_out_2_req_bits_addr),
    .io_out_2_req_bits_cmd(mmioXbar_io_out_2_req_bits_cmd),
    .io_out_2_req_bits_wmask(mmioXbar_io_out_2_req_bits_wmask),
    .io_out_2_req_bits_wdata(mmioXbar_io_out_2_req_bits_wdata),
    .io_out_2_resp_ready(mmioXbar_io_out_2_resp_ready),
    .io_out_2_resp_valid(mmioXbar_io_out_2_resp_valid),
    .io_out_2_resp_bits_cmd(mmioXbar_io_out_2_resp_bits_cmd),
    .io_out_2_resp_bits_rdata(mmioXbar_io_out_2_resp_bits_rdata)
  );
  AXI4CLINT clint ( // @[src/main/scala/system/NutShell.scala 113:21]
    .clock(clint_clock),
    .reset(clint_reset),
    .io__in_aw_ready(clint_io__in_aw_ready),
    .io__in_aw_valid(clint_io__in_aw_valid),
    .io__in_aw_bits_addr(clint_io__in_aw_bits_addr),
    .io__in_w_ready(clint_io__in_w_ready),
    .io__in_w_valid(clint_io__in_w_valid),
    .io__in_w_bits_data(clint_io__in_w_bits_data),
    .io__in_w_bits_strb(clint_io__in_w_bits_strb),
    .io__in_b_ready(clint_io__in_b_ready),
    .io__in_b_valid(clint_io__in_b_valid),
    .io__in_ar_ready(clint_io__in_ar_ready),
    .io__in_ar_valid(clint_io__in_ar_valid),
    .io__in_ar_bits_addr(clint_io__in_ar_bits_addr),
    .io__in_r_ready(clint_io__in_r_ready),
    .io__in_r_valid(clint_io__in_r_valid),
    .io__in_r_bits_data(clint_io__in_r_bits_data),
    .io__extra_mtip(clint_io__extra_mtip),
    .io__extra_msip(clint_io__extra_msip),
    .isWFI_0(clint_isWFI_0),
    .io_extra_mtip(clint_io_extra_mtip),
    .io_extra_msip(clint_io_extra_msip)
  );
  SimpleBus2AXI4Converter_1 clint_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(clint_io_in_bridge_clock),
    .reset(clint_io_in_bridge_reset),
    .io_in_req_ready(clint_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(clint_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(clint_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(clint_io_in_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(clint_io_in_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(clint_io_in_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(clint_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(clint_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(clint_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(clint_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(clint_io_in_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(clint_io_in_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(clint_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(clint_io_in_bridge_io_out_w_valid),
    .io_out_w_bits_data(clint_io_in_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(clint_io_in_bridge_io_out_w_bits_strb),
    .io_out_b_ready(clint_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(clint_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(clint_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(clint_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(clint_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(clint_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(clint_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(clint_io_in_bridge_io_out_r_bits_data)
  );
  AXI4PLIC plic ( // @[src/main/scala/system/NutShell.scala 120:20]
    .clock(plic_clock),
    .reset(plic_reset),
    .io__in_aw_ready(plic_io__in_aw_ready),
    .io__in_aw_valid(plic_io__in_aw_valid),
    .io__in_aw_bits_addr(plic_io__in_aw_bits_addr),
    .io__in_w_ready(plic_io__in_w_ready),
    .io__in_w_valid(plic_io__in_w_valid),
    .io__in_w_bits_data(plic_io__in_w_bits_data),
    .io__in_w_bits_strb(plic_io__in_w_bits_strb),
    .io__in_b_ready(plic_io__in_b_ready),
    .io__in_b_valid(plic_io__in_b_valid),
    .io__in_ar_ready(plic_io__in_ar_ready),
    .io__in_ar_valid(plic_io__in_ar_valid),
    .io__in_ar_bits_addr(plic_io__in_ar_bits_addr),
    .io__in_r_ready(plic_io__in_r_ready),
    .io__in_r_valid(plic_io__in_r_valid),
    .io__in_r_bits_data(plic_io__in_r_bits_data),
    .io__extra_meip_0(plic_io__extra_meip_0),
    .io_extra_meip_0(plic_io_extra_meip_0)
  );
  SimpleBus2AXI4Converter_2 plic_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(plic_io_in_bridge_clock),
    .reset(plic_io_in_bridge_reset),
    .io_in_req_ready(plic_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(plic_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(plic_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(plic_io_in_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(plic_io_in_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(plic_io_in_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(plic_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(plic_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(plic_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(plic_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(plic_io_in_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(plic_io_in_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(plic_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(plic_io_in_bridge_io_out_w_valid),
    .io_out_w_bits_data(plic_io_in_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(plic_io_in_bridge_io_out_w_bits_strb),
    .io_out_b_ready(plic_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(plic_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(plic_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(plic_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(plic_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(plic_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(plic_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(plic_io_in_bridge_io_out_r_bits_data)
  );
  assign io_mem_aw_valid = io_mem_bridge_io_out_aw_valid; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_aw_bits_addr = io_mem_bridge_io_out_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_w_valid = io_mem_bridge_io_out_w_valid; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_w_bits_data = io_mem_bridge_io_out_w_bits_data; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_w_bits_strb = io_mem_bridge_io_out_w_bits_strb; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_w_bits_last = io_mem_bridge_io_out_w_bits_last; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_ar_valid = io_mem_bridge_io_out_ar_valid; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_ar_bits_addr = io_mem_bridge_io_out_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_ar_bits_len = io_mem_bridge_io_out_ar_bits_len; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_ar_bits_size = io_mem_bridge_io_out_ar_bits_size; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mmio_req_valid = mmioXbar_io_out_2_req_valid; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_req_bits_addr = mmioXbar_io_out_2_req_bits_addr; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_req_bits_cmd = mmioXbar_io_out_2_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_req_bits_wmask = mmioXbar_io_out_2_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_req_bits_wdata = mmioXbar_io_out_2_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 111:18]
  assign io_mmio_resp_ready = mmioXbar_io_out_2_resp_ready; // @[src/main/scala/system/NutShell.scala 111:18]
  assign nutcore_clock = clock;
  assign nutcore_reset = reset;
  assign nutcore_io_imem_mem_req_ready = cohMg_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_valid = cohMg_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_bits_rdata = cohMg_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 56:15]
  assign nutcore_io_dmem_mem_req_ready = xbar_io_in_1_req_ready; // @[src/main/scala/system/NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_valid = xbar_io_in_1_resp_valid; // @[src/main/scala/system/NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_bits_cmd = xbar_io_in_1_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_bits_rdata = xbar_io_in_1_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 59:17]
  assign nutcore_io_mmio_req_ready = mmioXbar_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_valid = mmioXbar_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_bits_cmd = mmioXbar_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_bits_rdata = mmioXbar_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 107:18]
  assign nutcore_io_extra_meip_0 = plic_io_extra_meip_0;
  assign nutcore_io_extra_mtip = clint_io_extra_mtip;
  assign nutcore_io_extra_msip = clint_io_extra_msip;
  assign cohMg_clock = clock;
  assign cohMg_reset = reset;
  assign cohMg_io_in_req_valid = nutcore_io_imem_mem_req_valid; // @[src/main/scala/system/NutShell.scala 56:15]
  assign cohMg_io_in_req_bits_addr = nutcore_io_imem_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 56:15]
  assign cohMg_io_out_mem_req_ready = xbar_io_in_0_req_ready; // @[src/main/scala/system/NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_valid = xbar_io_in_0_resp_valid; // @[src/main/scala/system/NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_bits_cmd = xbar_io_in_0_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_bits_rdata = xbar_io_in_0_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 58:17]
  assign xbar_clock = clock;
  assign xbar_reset = reset;
  assign xbar_io_in_0_req_valid = cohMg_io_out_mem_req_valid; // @[src/main/scala/system/NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_addr = cohMg_io_out_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 58:17]
  assign xbar_io_in_1_req_valid = nutcore_io_dmem_mem_req_valid; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_addr = nutcore_io_dmem_mem_req_bits_addr; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_size = nutcore_io_dmem_mem_req_bits_size; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_cmd = nutcore_io_dmem_mem_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_wmask = nutcore_io_dmem_mem_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_wdata = nutcore_io_dmem_mem_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 59:17]
  assign xbar_io_out_req_ready = memAddrMap_io_in_req_ready; // @[src/main/scala/system/NutShell.scala 94:20]
  assign xbar_io_out_resp_valid = memAddrMap_io_in_resp_valid; // @[src/main/scala/system/NutShell.scala 94:20]
  assign xbar_io_out_resp_bits_cmd = memAddrMap_io_in_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 94:20]
  assign xbar_io_out_resp_bits_rdata = memAddrMap_io_in_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 94:20]
  assign axi2sb_clock = clock;
  assign axi2sb_reset = reset;
  assign memport_bridge_clock = clock;
  assign memport_bridge_reset = reset;
  assign memAddrMap_clock = clock;
  assign memAddrMap_reset = reset;
  assign memAddrMap_io_in_req_valid = xbar_io_out_req_valid; // @[src/main/scala/system/NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_addr = xbar_io_out_req_bits_addr; // @[src/main/scala/system/NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_size = xbar_io_out_req_bits_size; // @[src/main/scala/system/NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_cmd = xbar_io_out_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_wmask = xbar_io_out_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_wdata = xbar_io_out_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 94:20]
  assign memAddrMap_io_out_req_ready = io_mem_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_valid = io_mem_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_bits_cmd = io_mem_bridge_io_in_resp_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_bits_rdata = io_mem_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_clock = clock;
  assign io_mem_bridge_reset = reset;
  assign io_mem_bridge_io_in_req_valid = memAddrMap_io_out_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_in_req_bits_addr = memAddrMap_io_out_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_in_req_bits_size = memAddrMap_io_out_req_bits_size; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_in_req_bits_cmd = memAddrMap_io_out_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_in_req_bits_wmask = memAddrMap_io_out_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_in_req_bits_wdata = memAddrMap_io_out_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign io_mem_bridge_io_out_aw_ready = io_mem_aw_ready; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_w_ready = io_mem_w_ready; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_b_valid = io_mem_b_valid; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_r_valid = io_mem_r_valid; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_r_bits_data = io_mem_r_bits_data; // @[src/main/scala/system/NutShell.scala 95:10]
  assign io_mem_bridge_io_out_r_bits_last = io_mem_r_bits_last; // @[src/main/scala/system/NutShell.scala 95:10]
  assign mmioXbar_clock = clock;
  assign mmioXbar_reset = reset;
  assign mmioXbar_io_in_req_valid = nutcore_io_mmio_req_valid; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_addr = nutcore_io_mmio_req_bits_addr; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_cmd = nutcore_io_mmio_req_bits_cmd; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_wmask = nutcore_io_mmio_req_bits_wmask; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_wdata = nutcore_io_mmio_req_bits_wdata; // @[src/main/scala/system/NutShell.scala 107:18]
  assign mmioXbar_io_out_0_req_ready = clint_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_0_resp_valid = clint_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_0_resp_bits_rdata = clint_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_req_ready = plic_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_resp_valid = plic_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_resp_bits_rdata = plic_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign mmioXbar_io_out_2_req_ready = io_mmio_req_ready; // @[src/main/scala/system/NutShell.scala 111:18]
  assign mmioXbar_io_out_2_resp_valid = io_mmio_resp_valid; // @[src/main/scala/system/NutShell.scala 111:18]
  assign mmioXbar_io_out_2_resp_bits_cmd = io_mmio_resp_bits_cmd; // @[src/main/scala/system/NutShell.scala 111:18]
  assign mmioXbar_io_out_2_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[src/main/scala/system/NutShell.scala 111:18]
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_io__in_aw_valid = clint_io_in_bridge_io_out_aw_valid; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_aw_bits_addr = clint_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_w_valid = clint_io_in_bridge_io_out_w_valid; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_w_bits_data = clint_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_w_bits_strb = clint_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_b_ready = clint_io_in_bridge_io_out_b_ready; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_ar_valid = clint_io_in_bridge_io_out_ar_valid; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_ar_bits_addr = clint_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io__in_r_ready = clint_io_in_bridge_io_out_r_ready; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_isWFI_0 = nutcore_isWFI;
  assign clint_io_in_bridge_clock = clock;
  assign clint_io_in_bridge_reset = reset;
  assign clint_io_in_bridge_io_in_req_valid = mmioXbar_io_out_0_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_in_req_bits_addr = mmioXbar_io_out_0_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_in_req_bits_cmd = mmioXbar_io_out_0_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_in_req_bits_wmask = mmioXbar_io_out_0_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_in_req_bits_wdata = mmioXbar_io_out_0_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_in_resp_ready = mmioXbar_io_out_0_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign clint_io_in_bridge_io_out_aw_ready = clint_io__in_aw_ready; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io_in_bridge_io_out_w_ready = clint_io__in_w_ready; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io_in_bridge_io_out_b_valid = clint_io__in_b_valid; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io_in_bridge_io_out_ar_ready = clint_io__in_ar_ready; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io_in_bridge_io_out_r_valid = clint_io__in_r_valid; // @[src/main/scala/system/NutShell.scala 114:15]
  assign clint_io_in_bridge_io_out_r_bits_data = clint_io__in_r_bits_data; // @[src/main/scala/system/NutShell.scala 114:15]
  assign plic_clock = clock;
  assign plic_reset = reset;
  assign plic_io__in_aw_valid = plic_io_in_bridge_io_out_aw_valid; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_aw_bits_addr = plic_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_w_valid = plic_io_in_bridge_io_out_w_valid; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_w_bits_data = plic_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_w_bits_strb = plic_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_b_ready = plic_io_in_bridge_io_out_b_ready; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_ar_valid = plic_io_in_bridge_io_out_ar_valid; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_ar_bits_addr = plic_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io__in_r_ready = plic_io_in_bridge_io_out_r_ready; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_clock = clock;
  assign plic_io_in_bridge_reset = reset;
  assign plic_io_in_bridge_io_in_req_valid = mmioXbar_io_out_1_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_in_req_bits_addr = mmioXbar_io_out_1_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_in_req_bits_cmd = mmioXbar_io_out_1_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_in_req_bits_wmask = mmioXbar_io_out_1_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_in_req_bits_wdata = mmioXbar_io_out_1_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_in_resp_ready = mmioXbar_io_out_1_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign plic_io_in_bridge_io_out_aw_ready = plic_io__in_aw_ready; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_io_out_w_ready = plic_io__in_w_ready; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_io_out_b_valid = plic_io__in_b_valid; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_io_out_ar_ready = plic_io__in_ar_ready; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_io_out_r_valid = plic_io__in_r_valid; // @[src/main/scala/system/NutShell.scala 121:14]
  assign plic_io_in_bridge_io_out_r_bits_data = plic_io__in_r_bits_data; // @[src/main/scala/system/NutShell.scala 121:14]
endmodule
module DifftestMem1P(
  input         clock,
  input         reset,
  input         read_valid, // @[difftest/src/main/scala/common/Mem.scala 199:16]
  input  [63:0] read_index, // @[difftest/src/main/scala/common/Mem.scala 199:16]
  output [63:0] read_data_0, // @[difftest/src/main/scala/common/Mem.scala 199:16]
  input         write_valid, // @[difftest/src/main/scala/common/Mem.scala 204:17]
  input  [63:0] write_index, // @[difftest/src/main/scala/common/Mem.scala 204:17]
  input  [63:0] write_data_0, // @[difftest/src/main/scala/common/Mem.scala 204:17]
  input  [63:0] write_mask_0 // @[difftest/src/main/scala/common/Mem.scala 204:17]
);
  wire  helper_0_r_enable; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire [63:0] helper_0_r_index; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire [63:0] helper_0_r_data; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire  helper_0_w_enable; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire [63:0] helper_0_w_index; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire [63:0] helper_0_w_data; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire [63:0] helper_0_w_mask; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire  helper_0_clock; // @[difftest/src/main/scala/common/Mem.scala 197:49]
  wire  _T_1 = ~reset; // @[difftest/src/main/scala/common/Mem.scala 214:16]
  wire [64:0] _T_3 = read_index * 1'h1; // @[difftest/src/main/scala/common/Mem.scala 215:26]
  wire [65:0] _T_4 = {{1'd0}, _T_3}; // @[difftest/src/main/scala/common/Mem.scala 215:39]
  wire [64:0] _T_9 = write_index * 1'h1; // @[difftest/src/main/scala/common/Mem.scala 223:27]
  wire [65:0] _T_10 = {{1'd0}, _T_9}; // @[difftest/src/main/scala/common/Mem.scala 223:40]
  MemRWHelper helper_0 ( // @[difftest/src/main/scala/common/Mem.scala 197:49]
    .r_enable(helper_0_r_enable),
    .r_index(helper_0_r_index),
    .r_data(helper_0_r_data),
    .w_enable(helper_0_w_enable),
    .w_index(helper_0_w_index),
    .w_data(helper_0_w_data),
    .w_mask(helper_0_w_mask),
    .clock(helper_0_clock)
  );
  assign read_data_0 = helper_0_r_data; // @[difftest/src/main/scala/common/Mem.scala 211:13]
  assign helper_0_r_enable = ~reset & read_valid; // @[difftest/src/main/scala/common/Mem.scala 214:30]
  assign helper_0_r_index = _T_4[63:0]; // @[difftest/src/main/scala/common/Mem.scala 102:13]
  assign helper_0_w_enable = _T_1 & write_valid; // @[difftest/src/main/scala/common/Mem.scala 222:30]
  assign helper_0_w_index = _T_10[63:0]; // @[difftest/src/main/scala/common/Mem.scala 150:13]
  assign helper_0_w_data = write_data_0; // @[difftest/src/main/scala/common/Mem.scala 151:12]
  assign helper_0_w_mask = write_mask_0; // @[difftest/src/main/scala/common/Mem.scala 152:12]
  assign helper_0_clock = clock; // @[difftest/src/main/scala/common/Mem.scala 220:13]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1 & ~(~read_valid | ~write_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed: read and write come at the same cycle\n    at Mem.scala:263 assert(!read.valid || !write.valid, \"read and write come at the same cycle\")\n"
            ); // @[difftest/src/main/scala/common/Mem.scala 263:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge clock) begin
    //
    if (_T_1) begin
      assert(~read_valid | ~write_valid); // @[difftest/src/main/scala/common/Mem.scala 263:9]
    end
  end
endmodule
module AXI4RAM(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_bits_last, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_in_ar_bits_len, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [2:0]  io_in_ar_bits_size, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_bits_last // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
`endif // RANDOMIZE_REG_INIT
  wire  rdata_mem_clock; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire  rdata_mem_reset; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire  rdata_mem_read_valid; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire [63:0] rdata_mem_read_index; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire [63:0] rdata_mem_read_data_0; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire  rdata_mem_write_valid; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire [63:0] rdata_mem_write_index; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire [63:0] rdata_mem_write_data_0; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire [63:0] rdata_mem_write_mask_0; // @[difftest/src/main/scala/common/Mem.scala 322:36]
  wire [7:0] _fullMask_T_8 = io_in_w_bits_strb[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_9 = io_in_w_bits_strb[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_10 = io_in_w_bits_strb[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_11 = io_in_w_bits_strb[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_12 = io_in_w_bits_strb[4] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_13 = io_in_w_bits_strb[5] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_14 = io_in_w_bits_strb[6] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _fullMask_T_15 = io_in_w_bits_strb[7] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [31:0] fullMask_lo = {_fullMask_T_11,_fullMask_T_10,_fullMask_T_9,_fullMask_T_8}; // @[src/main/scala/utils/BitUtils.scala 27:27]
  wire [31:0] fullMask_hi = {_fullMask_T_15,_fullMask_T_14,_fullMask_T_13,_fullMask_T_12}; // @[src/main/scala/utils/BitUtils.scala 27:27]
  reg [7:0] c_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  reg [7:0] readBeatCnt; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  _len_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg [7:0] len_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [7:0] _GEN_0 = _len_T ? io_in_ar_bits_len : len_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  reg [1:0] burst_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [1:0] _GEN_1 = _len_T ? 2'h2 : burst_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  wire [31:0] _wrapAddr_WIRE = {{24'd0}, io_in_ar_bits_len}; // @[src/main/scala/device/AXI4Slave.scala 45:{69,69}]
  wire [38:0] _GEN_42 = {{7'd0}, _wrapAddr_WIRE}; // @[src/main/scala/device/AXI4Slave.scala 45:89]
  wire [38:0] _wrapAddr_T = _GEN_42 << io_in_ar_bits_size; // @[src/main/scala/device/AXI4Slave.scala 45:89]
  wire [38:0] _wrapAddr_T_1 = ~_wrapAddr_T; // @[src/main/scala/device/AXI4Slave.scala 45:42]
  wire [38:0] _GEN_34 = {{7'd0}, io_in_ar_bits_addr}; // @[src/main/scala/device/AXI4Slave.scala 45:40]
  wire [38:0] wrapAddr = _GEN_34 & _wrapAddr_T_1; // @[src/main/scala/device/AXI4Slave.scala 45:40]
  reg [38:0] raddr_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [38:0] _GEN_2 = _len_T ? wrapAddr : raddr_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  wire [7:0] _value_T_1 = readBeatCnt + 8'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [7:0] _GEN_3 = _GEN_1 == 2'h2 & readBeatCnt == _GEN_0 ? 8'h0 : _value_T_1; // @[src/main/scala/device/AXI4Slave.scala 50:{77,93} src/main/scala/chisel3/util/Counter.scala 77:15]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  ren = ren_REG | io_in_r_valid & ~io_in_r_bits_last; // @[src/main/scala/device/AXI4Slave.scala 73:46]
  wire [7:0] _GEN_4 = ren ? _GEN_3 : readBeatCnt; // @[src/main/scala/device/AXI4Slave.scala 48:18 src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [7:0] _value_T_3 = c_value + 8'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [31:0] _value_T_4 = io_in_ar_bits_addr >> io_in_ar_bits_size; // @[src/main/scala/device/AXI4Slave.scala 57:45]
  wire [31:0] _GEN_35 = {{24'd0}, io_in_ar_bits_len}; // @[src/main/scala/device/AXI4Slave.scala 57:67]
  wire [31:0] _value_T_5 = _value_T_4 & _GEN_35; // @[src/main/scala/device/AXI4Slave.scala 57:67]
  wire  _T_5 = io_in_ar_bits_len != 8'h0; // @[src/main/scala/device/AXI4Slave.scala 58:32]
  wire  _T_11 = io_in_ar_bits_len == 8'h7; // @[src/main/scala/device/AXI4Slave.scala 60:30]
  wire  _T_12 = io_in_ar_bits_len == 8'h1 | io_in_ar_bits_len == 8'h3 | _T_11; // @[src/main/scala/device/AXI4Slave.scala 59:71]
  wire  _T_14 = _T_12 | io_in_ar_bits_len == 8'hf; // @[src/main/scala/device/AXI4Slave.scala 60:38]
  wire [31:0] _GEN_7 = _len_T ? _value_T_5 : {{24'd0}, _GEN_4}; // @[src/main/scala/device/AXI4Slave.scala 56:29 57:23]
  wire  _r_busy_T_2 = io_in_r_valid & io_in_r_bits_last; // @[src/main/scala/device/AXI4Slave.scala 70:56]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_8 = _r_busy_T_2 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_9 = _len_T | _GEN_8; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_r_valid_T_2 = ren & (_len_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_10 = io_in_r_valid ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_11 = _io_in_r_valid_T_2 | _GEN_10; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [7:0] writeBeatCnt; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  _waddr_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg [31:0] waddr_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [31:0] _GEN_12 = _waddr_T ? io_in_aw_bits_addr : waddr_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  wire  _T_18 = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [7:0] _value_T_7 = writeBeatCnt + 8'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_15 = io_in_b_valid ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_16 = _waddr_T | _GEN_15; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T_1 = _T_18 & io_in_w_bits_last; // @[src/main/scala/device/AXI4Slave.scala 97:43]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_17 = io_in_b_valid ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_18 = _io_in_b_valid_T_1 | _GEN_17; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire [31:0] _wIdx_T = _GEN_12 & 32'h7fffffff; // @[src/main/scala/device/AXI4RAM.scala 32:33]
  wire [28:0] _GEN_36 = {{21'd0}, writeBeatCnt}; // @[src/main/scala/device/AXI4RAM.scala 35:27]
  wire [28:0] wIdx = _wIdx_T[31:3] + _GEN_36; // @[src/main/scala/device/AXI4RAM.scala 35:27]
  wire [38:0] _rIdx_T = _GEN_2 & 39'h7fffffff; // @[src/main/scala/device/AXI4RAM.scala 32:33]
  wire [35:0] _GEN_37 = {{28'd0}, readBeatCnt}; // @[src/main/scala/device/AXI4RAM.scala 36:27]
  wire [35:0] rIdx = _rIdx_T[38:3] + _GEN_37; // @[src/main/scala/device/AXI4RAM.scala 36:27]
  wire  _wen_T_1 = wIdx < 29'h10000000; // @[src/main/scala/device/AXI4RAM.scala 33:32]
  wire [31:0] rdata_lo = {io_in_w_bits_data[31:24],io_in_w_bits_data[23:16],io_in_w_bits_data[15:8],io_in_w_bits_data[7:
    0]}; // @[difftest/src/main/scala/common/Mem.scala 244:41]
  wire [31:0] rdata_hi = {io_in_w_bits_data[63:56],io_in_w_bits_data[55:48],io_in_w_bits_data[47:40],io_in_w_bits_data[
    39:32]}; // @[difftest/src/main/scala/common/Mem.scala 244:41]
  reg  rdata_REG; // @[difftest/src/main/scala/common/Mem.scala 238:16]
  reg  rdata_REG_1; // @[difftest/src/main/scala/common/Mem.scala 238:61]
  reg [63:0] rdata_r_0; // @[difftest/src/main/scala/common/Mem.scala 238:42]
  wire [63:0] _rdata_T_28_0 = rdata_REG ? rdata_mem_read_data_0 : rdata_r_0; // @[difftest/src/main/scala/common/Mem.scala 238:8]
  wire [31:0] rdata_lo_2 = {_rdata_T_28_0[31:24],_rdata_T_28_0[23:16],_rdata_T_28_0[15:8],_rdata_T_28_0[7:0]}; // @[src/main/scala/device/AXI4RAM.scala 48:32]
  wire [31:0] rdata_hi_2 = {_rdata_T_28_0[63:56],_rdata_T_28_0[55:48],_rdata_T_28_0[47:40],_rdata_T_28_0[39:32]}; // @[src/main/scala/device/AXI4RAM.scala 48:32]
  wire [31:0] _GEN_38 = reset ? 32'h0 : _GEN_7; // @[src/main/scala/chisel3/util/Counter.scala 61:{40,40}]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [7:0] c_value_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [7:0] c_value_t = c_value ^ c_value_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  toggle_10635_clock;
  wire  toggle_10635_reset;
  wire [7:0] toggle_10635_valid;
  reg [7:0] toggle_10635_valid_reg;
  reg [7:0] readBeatCnt_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [7:0] readBeatCnt_t = readBeatCnt ^ readBeatCnt_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  toggle_10643_clock;
  wire  toggle_10643_reset;
  wire [7:0] toggle_10643_valid;
  reg [7:0] toggle_10643_valid_reg;
  reg [7:0] len_r_p; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [7:0] len_r_t = len_r ^ len_r_p; // @[src/main/scala/utils/Hold.scala 23:65]
  wire  toggle_10651_clock;
  wire  toggle_10651_reset;
  wire [7:0] toggle_10651_valid;
  reg [7:0] toggle_10651_valid_reg;
  reg [1:0] burst_r_p; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [1:0] burst_r_t = burst_r ^ burst_r_p; // @[src/main/scala/utils/Hold.scala 23:65]
  wire  toggle_10659_clock;
  wire  toggle_10659_reset;
  wire [1:0] toggle_10659_valid;
  reg [1:0] toggle_10659_valid_reg;
  reg [38:0] raddr_r_p; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [38:0] raddr_r_t = raddr_r ^ raddr_r_p; // @[src/main/scala/utils/Hold.scala 23:65]
  wire  toggle_10661_clock;
  wire  toggle_10661_reset;
  wire [38:0] toggle_10661_valid;
  reg [38:0] toggle_10661_valid_reg;
  reg  ren_REG_p; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  ren_REG_t = ren_REG ^ ren_REG_p; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  toggle_10700_clock;
  wire  toggle_10700_reset;
  wire  toggle_10700_valid;
  reg  toggle_10700_valid_reg;
  reg  r_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  r_busy_t = r_busy ^ r_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10701_clock;
  wire  toggle_10701_reset;
  wire  toggle_10701_valid;
  reg  toggle_10701_valid_reg;
  reg  io_in_r_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  io_in_r_valid_r_t = io_in_r_valid_r ^ io_in_r_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10702_clock;
  wire  toggle_10702_reset;
  wire  toggle_10702_valid;
  reg  toggle_10702_valid_reg;
  reg [7:0] writeBeatCnt_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [7:0] writeBeatCnt_t = writeBeatCnt ^ writeBeatCnt_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  toggle_10703_clock;
  wire  toggle_10703_reset;
  wire [7:0] toggle_10703_valid;
  reg [7:0] toggle_10703_valid_reg;
  reg [31:0] waddr_r_p; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [31:0] waddr_r_t = waddr_r ^ waddr_r_p; // @[src/main/scala/utils/Hold.scala 23:65]
  wire  toggle_10711_clock;
  wire  toggle_10711_reset;
  wire [31:0] toggle_10711_valid;
  reg [31:0] toggle_10711_valid_reg;
  reg  w_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  w_busy_t = w_busy ^ w_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10743_clock;
  wire  toggle_10743_reset;
  wire  toggle_10743_valid;
  reg  toggle_10743_valid_reg;
  reg  io_in_b_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  io_in_b_valid_r_t = io_in_b_valid_r ^ io_in_b_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10744_clock;
  wire  toggle_10744_reset;
  wire  toggle_10744_valid;
  reg  toggle_10744_valid_reg;
  reg  rdata_REG_p; // @[difftest/src/main/scala/common/Mem.scala 238:16]
  wire  rdata_REG_t = rdata_REG ^ rdata_REG_p; // @[difftest/src/main/scala/common/Mem.scala 238:16]
  wire  toggle_10745_clock;
  wire  toggle_10745_reset;
  wire  toggle_10745_valid;
  reg  toggle_10745_valid_reg;
  reg  rdata_REG_1_p; // @[difftest/src/main/scala/common/Mem.scala 238:61]
  wire  rdata_REG_1_t = rdata_REG_1 ^ rdata_REG_1_p; // @[difftest/src/main/scala/common/Mem.scala 238:61]
  wire  toggle_10746_clock;
  wire  toggle_10746_reset;
  wire  toggle_10746_valid;
  reg  toggle_10746_valid_reg;
  reg [63:0] rdata_r_0_p; // @[difftest/src/main/scala/common/Mem.scala 238:42]
  wire [63:0] rdata_r_0_t = rdata_r_0 ^ rdata_r_0_p; // @[difftest/src/main/scala/common/Mem.scala 238:42]
  wire  toggle_10747_clock;
  wire  toggle_10747_reset;
  wire [63:0] toggle_10747_valid;
  reg [63:0] toggle_10747_valid_reg;
  DifftestMem1P rdata_mem ( // @[difftest/src/main/scala/common/Mem.scala 322:36]
    .clock(rdata_mem_clock),
    .reset(rdata_mem_reset),
    .read_valid(rdata_mem_read_valid),
    .read_index(rdata_mem_read_index),
    .read_data_0(rdata_mem_read_data_0),
    .write_valid(rdata_mem_write_valid),
    .write_index(rdata_mem_write_index),
    .write_data_0(rdata_mem_write_data_0),
    .write_mask_0(rdata_mem_write_mask_0)
  );
  GEN_w8_toggle #(.COVER_INDEX(10635)) toggle_10635 (
    .clock(toggle_10635_clock),
    .reset(toggle_10635_reset),
    .valid(toggle_10635_valid)
  );
  GEN_w8_toggle #(.COVER_INDEX(10643)) toggle_10643 (
    .clock(toggle_10643_clock),
    .reset(toggle_10643_reset),
    .valid(toggle_10643_valid)
  );
  GEN_w8_toggle #(.COVER_INDEX(10651)) toggle_10651 (
    .clock(toggle_10651_clock),
    .reset(toggle_10651_reset),
    .valid(toggle_10651_valid)
  );
  GEN_w2_toggle #(.COVER_INDEX(10659)) toggle_10659 (
    .clock(toggle_10659_clock),
    .reset(toggle_10659_reset),
    .valid(toggle_10659_valid)
  );
  GEN_w39_toggle #(.COVER_INDEX(10661)) toggle_10661 (
    .clock(toggle_10661_clock),
    .reset(toggle_10661_reset),
    .valid(toggle_10661_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10700)) toggle_10700 (
    .clock(toggle_10700_clock),
    .reset(toggle_10700_reset),
    .valid(toggle_10700_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10701)) toggle_10701 (
    .clock(toggle_10701_clock),
    .reset(toggle_10701_reset),
    .valid(toggle_10701_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10702)) toggle_10702 (
    .clock(toggle_10702_clock),
    .reset(toggle_10702_reset),
    .valid(toggle_10702_valid)
  );
  GEN_w8_toggle #(.COVER_INDEX(10703)) toggle_10703 (
    .clock(toggle_10703_clock),
    .reset(toggle_10703_reset),
    .valid(toggle_10703_valid)
  );
  GEN_w32_toggle #(.COVER_INDEX(10711)) toggle_10711 (
    .clock(toggle_10711_clock),
    .reset(toggle_10711_reset),
    .valid(toggle_10711_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10743)) toggle_10743 (
    .clock(toggle_10743_clock),
    .reset(toggle_10743_reset),
    .valid(toggle_10743_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10744)) toggle_10744 (
    .clock(toggle_10744_clock),
    .reset(toggle_10744_reset),
    .valid(toggle_10744_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10745)) toggle_10745 (
    .clock(toggle_10745_clock),
    .reset(toggle_10745_reset),
    .valid(toggle_10745_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10746)) toggle_10746 (
    .clock(toggle_10746_clock),
    .reset(toggle_10746_reset),
    .valid(toggle_10746_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(10747)) toggle_10747 (
    .clock(toggle_10747_clock),
    .reset(toggle_10747_reset),
    .valid(toggle_10747_valid)
  );
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = 1'h1; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = {rdata_hi_2,rdata_lo_2}; // @[src/main/scala/device/AXI4RAM.scala 48:32]
  assign io_in_r_bits_last = c_value == _GEN_0; // @[src/main/scala/device/AXI4Slave.scala 47:36]
  assign rdata_mem_clock = clock;
  assign rdata_mem_reset = reset;
  assign rdata_mem_read_valid = ren_REG | io_in_r_valid & ~io_in_r_bits_last; // @[src/main/scala/device/AXI4Slave.scala 73:46]
  assign rdata_mem_read_index = {{28'd0}, rIdx}; // @[difftest/src/main/scala/common/Mem.scala 237:16]
  assign rdata_mem_write_valid = _T_18 & _wen_T_1; // @[src/main/scala/device/AXI4RAM.scala 37:25]
  assign rdata_mem_write_index = {{35'd0}, wIdx};
  assign rdata_mem_write_data_0 = {rdata_hi,rdata_lo}; // @[difftest/src/main/scala/common/Mem.scala 244:41]
  assign rdata_mem_write_mask_0 = {fullMask_hi,fullMask_lo}; // @[difftest/src/main/scala/common/Mem.scala 248:65]
  assign toggle_10635_clock = clock;
  assign toggle_10635_reset = reset;
  assign toggle_10635_valid = c_value ^ toggle_10635_valid_reg;
  assign toggle_10643_clock = clock;
  assign toggle_10643_reset = reset;
  assign toggle_10643_valid = readBeatCnt ^ toggle_10643_valid_reg;
  assign toggle_10651_clock = clock;
  assign toggle_10651_reset = reset;
  assign toggle_10651_valid = len_r ^ toggle_10651_valid_reg;
  assign toggle_10659_clock = clock;
  assign toggle_10659_reset = reset;
  assign toggle_10659_valid = burst_r ^ toggle_10659_valid_reg;
  assign toggle_10661_clock = clock;
  assign toggle_10661_reset = reset;
  assign toggle_10661_valid = raddr_r ^ toggle_10661_valid_reg;
  assign toggle_10700_clock = clock;
  assign toggle_10700_reset = reset;
  assign toggle_10700_valid = ren_REG ^ toggle_10700_valid_reg;
  assign toggle_10701_clock = clock;
  assign toggle_10701_reset = reset;
  assign toggle_10701_valid = r_busy ^ toggle_10701_valid_reg;
  assign toggle_10702_clock = clock;
  assign toggle_10702_reset = reset;
  assign toggle_10702_valid = io_in_r_valid_r ^ toggle_10702_valid_reg;
  assign toggle_10703_clock = clock;
  assign toggle_10703_reset = reset;
  assign toggle_10703_valid = writeBeatCnt ^ toggle_10703_valid_reg;
  assign toggle_10711_clock = clock;
  assign toggle_10711_reset = reset;
  assign toggle_10711_valid = waddr_r ^ toggle_10711_valid_reg;
  assign toggle_10743_clock = clock;
  assign toggle_10743_reset = reset;
  assign toggle_10743_valid = w_busy ^ toggle_10743_valid_reg;
  assign toggle_10744_clock = clock;
  assign toggle_10744_reset = reset;
  assign toggle_10744_valid = io_in_b_valid_r ^ toggle_10744_valid_reg;
  assign toggle_10745_clock = clock;
  assign toggle_10745_reset = reset;
  assign toggle_10745_valid = rdata_REG ^ toggle_10745_valid_reg;
  assign toggle_10746_clock = clock;
  assign toggle_10746_reset = reset;
  assign toggle_10746_valid = rdata_REG_1 ^ toggle_10746_valid_reg;
  assign toggle_10747_clock = clock;
  assign toggle_10747_reset = reset;
  assign toggle_10747_valid = rdata_r_0 ^ toggle_10747_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      c_value <= 8'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (io_in_r_valid) begin // @[src/main/scala/device/AXI4Slave.scala 52:28]
      if (io_in_r_bits_last) begin // @[src/main/scala/device/AXI4Slave.scala 54:33]
        c_value <= 8'h0; // @[src/main/scala/device/AXI4Slave.scala 54:43]
      end else begin
        c_value <= _value_T_3; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
      end
    end
    readBeatCnt <= _GEN_38[7:0]; // @[src/main/scala/chisel3/util/Counter.scala 61:{40,40}]
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      len_r <= 8'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_len_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      len_r <= io_in_ar_bits_len; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      burst_r <= 2'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_len_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      burst_r <= 2'h2; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      raddr_r <= 39'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_len_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      raddr_r <= wrapAddr; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _len_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_9;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_11;
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      writeBeatCnt <= 8'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_T_18) begin // @[src/main/scala/device/AXI4Slave.scala 82:28]
      if (io_in_w_bits_last) begin // @[src/main/scala/device/AXI4Slave.scala 84:33]
        writeBeatCnt <= 8'h0; // @[src/main/scala/device/AXI4Slave.scala 84:43]
      end else begin
        writeBeatCnt <= _value_T_7; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
      end
    end
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      waddr_r <= 32'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_waddr_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      waddr_r <= io_in_aw_bits_addr; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_16;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_18;
    end
    rdata_REG <= ren_REG | io_in_r_valid & ~io_in_r_bits_last; // @[src/main/scala/device/AXI4Slave.scala 73:46]
    rdata_REG_1 <= ren_REG | io_in_r_valid & ~io_in_r_bits_last; // @[src/main/scala/device/AXI4Slave.scala 73:46]
    if (rdata_REG_1) begin // @[difftest/src/main/scala/common/Mem.scala 238:42]
      rdata_r_0 <= rdata_mem_read_data_0; // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_len_T & _T_5 & ~reset & ~_T_14) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at AXI4Slave.scala:59 assert(axi4.ar.bits.len === 1.U || axi4.ar.bits.len === 3.U ||\n"
            ); // @[src/main/scala/device/AXI4Slave.scala 59:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    c_value_p <= c_value; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    toggle_10635_valid_reg <= c_value;
    readBeatCnt_p <= readBeatCnt; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    toggle_10643_valid_reg <= readBeatCnt;
    len_r_p <= len_r; // @[src/main/scala/utils/Hold.scala 23:65]
    toggle_10651_valid_reg <= len_r;
    burst_r_p <= burst_r; // @[src/main/scala/utils/Hold.scala 23:65]
    toggle_10659_valid_reg <= burst_r;
    raddr_r_p <= raddr_r; // @[src/main/scala/utils/Hold.scala 23:65]
    toggle_10661_valid_reg <= raddr_r;
    ren_REG_p <= ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    toggle_10700_valid_reg <= ren_REG;
    r_busy_p <= r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10701_valid_reg <= r_busy;
    io_in_r_valid_r_p <= io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10702_valid_reg <= io_in_r_valid_r;
    writeBeatCnt_p <= writeBeatCnt; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    toggle_10703_valid_reg <= writeBeatCnt;
    waddr_r_p <= waddr_r; // @[src/main/scala/utils/Hold.scala 23:65]
    toggle_10711_valid_reg <= waddr_r;
    w_busy_p <= w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10743_valid_reg <= w_busy;
    io_in_b_valid_r_p <= io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10744_valid_reg <= io_in_b_valid_r;
    rdata_REG_p <= rdata_REG; // @[difftest/src/main/scala/common/Mem.scala 238:16]
    toggle_10745_valid_reg <= rdata_REG;
    rdata_REG_1_p <= rdata_REG_1; // @[difftest/src/main/scala/common/Mem.scala 238:61]
    toggle_10746_valid_reg <= rdata_REG_1;
    rdata_r_0_p <= rdata_r_0; // @[difftest/src/main/scala/common/Mem.scala 238:42]
    toggle_10747_valid_reg <= rdata_r_0;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  c_value = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  readBeatCnt = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  len_r = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  burst_r = _RAND_3[1:0];
  _RAND_4 = {2{`RANDOM}};
  raddr_r = _RAND_4[38:0];
  _RAND_5 = {1{`RANDOM}};
  ren_REG = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r_busy = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  writeBeatCnt = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  waddr_r = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  w_busy = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  rdata_REG = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  rdata_REG_1 = _RAND_13[0:0];
  _RAND_14 = {2{`RANDOM}};
  rdata_r_0 = _RAND_14[63:0];
  _RAND_15 = {1{`RANDOM}};
  c_value_p = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  toggle_10635_valid_reg = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  readBeatCnt_p = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  toggle_10643_valid_reg = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  len_r_p = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  toggle_10651_valid_reg = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  burst_r_p = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  toggle_10659_valid_reg = _RAND_22[1:0];
  _RAND_23 = {2{`RANDOM}};
  raddr_r_p = _RAND_23[38:0];
  _RAND_24 = {2{`RANDOM}};
  toggle_10661_valid_reg = _RAND_24[38:0];
  _RAND_25 = {1{`RANDOM}};
  ren_REG_p = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  toggle_10700_valid_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  r_busy_p = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  toggle_10701_valid_reg = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  io_in_r_valid_r_p = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  toggle_10702_valid_reg = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  writeBeatCnt_p = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  toggle_10703_valid_reg = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  waddr_r_p = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  toggle_10711_valid_reg = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  w_busy_p = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  toggle_10743_valid_reg = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  io_in_b_valid_r_p = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  toggle_10744_valid_reg = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  rdata_REG_p = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  toggle_10745_valid_reg = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  rdata_REG_1_p = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  toggle_10746_valid_reg = _RAND_42[0:0];
  _RAND_43 = {2{`RANDOM}};
  rdata_r_0_p = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  toggle_10747_valid_reg = _RAND_44[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_len_T & _T_5 & ~reset) begin
      assert(_T_14); // @[src/main/scala/device/AXI4Slave.scala 59:17]
    end
    //
    if (enToggle_past) begin
      cover(c_value_t[0]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(c_value_t[1]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(c_value_t[2]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(c_value_t[3]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(c_value_t[4]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(c_value_t[5]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(c_value_t[6]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(c_value_t[7]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(readBeatCnt_t[0]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(readBeatCnt_t[1]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(readBeatCnt_t[2]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(readBeatCnt_t[3]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(readBeatCnt_t[4]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(readBeatCnt_t[5]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(readBeatCnt_t[6]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(readBeatCnt_t[7]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(len_r_t[0]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(len_r_t[1]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(len_r_t[2]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(len_r_t[3]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(len_r_t[4]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(len_r_t[5]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(len_r_t[6]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(len_r_t[7]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(burst_r_t[0]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(burst_r_t[1]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[0]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[1]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[2]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[3]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[4]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[5]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[6]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[7]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[8]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[9]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[10]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[11]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[12]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[13]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[14]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[15]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[16]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[17]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[18]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[19]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[20]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[21]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[22]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[23]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[24]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[25]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[26]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[27]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[28]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[29]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[30]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[31]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[32]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[33]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[34]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[35]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[36]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[37]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(raddr_r_t[38]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(ren_REG_t); // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    //
    if (enToggle_past) begin
      cover(r_busy_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_valid_r_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(writeBeatCnt_t[0]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(writeBeatCnt_t[1]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(writeBeatCnt_t[2]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(writeBeatCnt_t[3]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(writeBeatCnt_t[4]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(writeBeatCnt_t[5]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(writeBeatCnt_t[6]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(writeBeatCnt_t[7]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[0]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[1]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[2]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[3]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[4]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[5]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[6]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[7]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[8]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[9]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[10]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[11]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[12]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[13]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[14]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[15]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[16]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[17]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[18]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[19]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[20]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[21]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[22]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[23]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[24]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[25]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[26]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[27]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[28]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[29]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[30]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(waddr_r_t[31]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(w_busy_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(io_in_b_valid_r_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(rdata_REG_t); // @[difftest/src/main/scala/common/Mem.scala 238:16]
    end
    //
    if (enToggle_past) begin
      cover(rdata_REG_1_t); // @[difftest/src/main/scala/common/Mem.scala 238:61]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[0]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[1]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[2]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[3]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[4]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[5]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[6]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[7]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[8]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[9]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[10]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[11]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[12]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[13]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[14]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[15]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[16]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[17]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[18]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[19]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[20]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[21]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[22]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[23]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[24]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[25]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[26]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[27]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[28]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[29]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[30]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[31]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[32]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[33]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[34]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[35]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[36]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[37]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[38]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[39]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[40]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[41]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[42]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[43]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[44]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[45]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[46]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[47]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[48]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[49]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[50]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[51]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[52]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[53]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[54]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[55]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[56]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[57]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[58]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[59]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[60]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[61]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[62]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
    //
    if (enToggle_past) begin
      cover(rdata_r_0_t[63]); // @[difftest/src/main/scala/common/Mem.scala 238:42]
    end
  end
endmodule
module LatencyPipe(
  input         clock,
  input         reset,
  input         io_in_valid, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input  [31:0] io_in_bits_addr, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input  [7:0]  io_in_bits_len, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input  [2:0]  io_in_bits_size, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output        io_out_valid, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output [31:0] io_out_bits_addr, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output [7:0]  io_out_bits_len, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output [2:0]  io_out_bits_size // @[src/main/scala/utils/LatencyPipe.scala 9:14]
);
  assign io_out_valid = io_in_valid; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  assign io_out_bits_addr = io_in_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  assign io_out_bits_len = io_in_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  assign io_out_bits_size = io_in_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
endmodule
module LatencyPipe_1(
  input         clock,
  input         reset,
  output        io_in_ready, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input         io_in_valid, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input  [31:0] io_in_bits_addr, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  input         io_out_ready, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output        io_out_valid, // @[src/main/scala/utils/LatencyPipe.scala 9:14]
  output [31:0] io_out_bits_addr // @[src/main/scala/utils/LatencyPipe.scala 9:14]
);
  assign io_in_ready = io_out_ready; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  assign io_out_valid = io_in_valid; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
  assign io_out_bits_addr = io_in_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 17:10]
endmodule
module AXI4Delayer(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_in_aw_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_in_w_ready, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_in_w_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [7:0]  io_in_w_bits_strb, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_in_w_bits_last, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_in_b_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_in_ar_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [7:0]  io_in_ar_bits_len, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [2:0]  io_in_ar_bits_size, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_in_r_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [63:0] io_in_r_bits_data, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_in_r_bits_last, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [31:0] io_out_aw_bits_addr, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_out_w_ready, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_out_w_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [63:0] io_out_w_bits_data, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [7:0]  io_out_w_bits_strb, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_out_w_bits_last, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_out_b_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [7:0]  io_out_ar_bits_len, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  output [2:0]  io_out_ar_bits_size, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_out_r_valid, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input  [63:0] io_out_r_bits_data, // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
  input         io_out_r_bits_last // @[src/main/scala/bus/axi4/Delayer.scala 10:14]
);
  wire  io_out_ar_pipe_clock; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_ar_pipe_reset; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_ar_pipe_io_in_valid; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [31:0] io_out_ar_pipe_io_in_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [7:0] io_out_ar_pipe_io_in_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [2:0] io_out_ar_pipe_io_in_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_ar_pipe_io_out_valid; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [31:0] io_out_ar_pipe_io_out_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [7:0] io_out_ar_pipe_io_out_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [2:0] io_out_ar_pipe_io_out_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_aw_pipe_clock; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_aw_pipe_reset; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_aw_pipe_io_in_ready; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_aw_pipe_io_in_valid; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [31:0] io_out_aw_pipe_io_in_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_aw_pipe_io_out_ready; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire  io_out_aw_pipe_io_out_valid; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  wire [31:0] io_out_aw_pipe_io_out_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 22:22]
  LatencyPipe io_out_ar_pipe ( // @[src/main/scala/utils/LatencyPipe.scala 22:22]
    .clock(io_out_ar_pipe_clock),
    .reset(io_out_ar_pipe_reset),
    .io_in_valid(io_out_ar_pipe_io_in_valid),
    .io_in_bits_addr(io_out_ar_pipe_io_in_bits_addr),
    .io_in_bits_len(io_out_ar_pipe_io_in_bits_len),
    .io_in_bits_size(io_out_ar_pipe_io_in_bits_size),
    .io_out_valid(io_out_ar_pipe_io_out_valid),
    .io_out_bits_addr(io_out_ar_pipe_io_out_bits_addr),
    .io_out_bits_len(io_out_ar_pipe_io_out_bits_len),
    .io_out_bits_size(io_out_ar_pipe_io_out_bits_size)
  );
  LatencyPipe_1 io_out_aw_pipe ( // @[src/main/scala/utils/LatencyPipe.scala 22:22]
    .clock(io_out_aw_pipe_clock),
    .reset(io_out_aw_pipe_reset),
    .io_in_ready(io_out_aw_pipe_io_in_ready),
    .io_in_valid(io_out_aw_pipe_io_in_valid),
    .io_in_bits_addr(io_out_aw_pipe_io_in_bits_addr),
    .io_out_ready(io_out_aw_pipe_io_out_ready),
    .io_out_valid(io_out_aw_pipe_io_out_valid),
    .io_out_bits_addr(io_out_aw_pipe_io_out_bits_addr)
  );
  assign io_in_aw_ready = io_out_aw_pipe_io_in_ready; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_in_w_ready = io_out_w_ready; // @[src/main/scala/bus/axi4/Delayer.scala 17:13]
  assign io_in_b_valid = io_out_b_valid; // @[src/main/scala/bus/axi4/Delayer.scala 18:13]
  assign io_in_r_valid = io_out_r_valid; // @[src/main/scala/bus/axi4/Delayer.scala 19:13]
  assign io_in_r_bits_data = io_out_r_bits_data; // @[src/main/scala/bus/axi4/Delayer.scala 19:13]
  assign io_in_r_bits_last = io_out_r_bits_last; // @[src/main/scala/bus/axi4/Delayer.scala 19:13]
  assign io_out_aw_valid = io_out_aw_pipe_io_out_valid; // @[src/main/scala/bus/axi4/Delayer.scala 16:13]
  assign io_out_aw_bits_addr = io_out_aw_pipe_io_out_bits_addr; // @[src/main/scala/bus/axi4/Delayer.scala 16:13]
  assign io_out_w_valid = io_in_w_valid; // @[src/main/scala/bus/axi4/Delayer.scala 17:13]
  assign io_out_w_bits_data = io_in_w_bits_data; // @[src/main/scala/bus/axi4/Delayer.scala 17:13]
  assign io_out_w_bits_strb = io_in_w_bits_strb; // @[src/main/scala/bus/axi4/Delayer.scala 17:13]
  assign io_out_w_bits_last = io_in_w_bits_last; // @[src/main/scala/bus/axi4/Delayer.scala 17:13]
  assign io_out_ar_valid = io_out_ar_pipe_io_out_valid; // @[src/main/scala/bus/axi4/Delayer.scala 15:13]
  assign io_out_ar_bits_addr = io_out_ar_pipe_io_out_bits_addr; // @[src/main/scala/bus/axi4/Delayer.scala 15:13]
  assign io_out_ar_bits_len = io_out_ar_pipe_io_out_bits_len; // @[src/main/scala/bus/axi4/Delayer.scala 15:13]
  assign io_out_ar_bits_size = io_out_ar_pipe_io_out_bits_size; // @[src/main/scala/bus/axi4/Delayer.scala 15:13]
  assign io_out_ar_pipe_clock = clock;
  assign io_out_ar_pipe_reset = reset;
  assign io_out_ar_pipe_io_in_valid = io_in_ar_valid; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_ar_pipe_io_in_bits_addr = io_in_ar_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_ar_pipe_io_in_bits_len = io_in_ar_bits_len; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_ar_pipe_io_in_bits_size = io_in_ar_bits_size; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_aw_pipe_clock = clock;
  assign io_out_aw_pipe_reset = reset;
  assign io_out_aw_pipe_io_in_valid = io_in_aw_valid; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_aw_pipe_io_in_bits_addr = io_in_aw_bits_addr; // @[src/main/scala/utils/LatencyPipe.scala 23:16]
  assign io_out_aw_pipe_io_out_ready = io_out_aw_ready; // @[src/main/scala/bus/axi4/Delayer.scala 16:13]
endmodule
module SimpleBusCrossbar1toN_1(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_in_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_in_resp_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_0_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_0_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_0_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_0_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_0_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_0_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_0_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_0_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_0_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_1_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_1_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_1_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_1_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_1_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_1_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_1_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_1_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_2_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_2_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_2_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_2_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_2_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_2_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_2_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_3_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_3_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_3_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_3_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_3_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_3_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_3_resp_bits_rdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_4_req_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_4_req_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [31:0] io_out_4_req_bits_addr, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [3:0]  io_out_4_req_bits_cmd, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [7:0]  io_out_4_req_bits_wmask, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output [63:0] io_out_4_req_bits_wdata, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  output        io_out_4_resp_ready, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input         io_out_4_resp_valid, // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
  input  [63:0] io_out_4_resp_bits_rdata // @[src/main/scala/bus/simplebus/Crossbar.scala 26:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
  wire  outMatchVec_0 = io_in_req_bits_addr >= 32'h40600000 & io_in_req_bits_addr < 32'h40600010; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_1 = io_in_req_bits_addr >= 32'h50000000 & io_in_req_bits_addr < 32'h50400000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_2 = io_in_req_bits_addr >= 32'h40001000 & io_in_req_bits_addr < 32'h40001008; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_3 = io_in_req_bits_addr >= 32'h40000000 & io_in_req_bits_addr < 32'h40001000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire  outMatchVec_4 = io_in_req_bits_addr >= 32'h40002000 & io_in_req_bits_addr < 32'h40003000; // @[src/main/scala/bus/simplebus/Crossbar.scala 37:34]
  wire [4:0] _outSelVec_enc_T = outMatchVec_4 ? 5'h10 : 5'h0; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _outSelVec_enc_T_1 = outMatchVec_3 ? 5'h8 : _outSelVec_enc_T; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _outSelVec_enc_T_2 = outMatchVec_2 ? 5'h4 : _outSelVec_enc_T_1; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _outSelVec_enc_T_3 = outMatchVec_1 ? 5'h2 : _outSelVec_enc_T_2; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] outSelVec_enc = outMatchVec_0 ? 5'h1 : _outSelVec_enc_T_3; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire  outSelVec_0 = outSelVec_enc[0]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_1 = outSelVec_enc[1]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_2 = outSelVec_enc[2]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_3 = outSelVec_enc[3]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  outSelVec_4 = outSelVec_enc[4]; // @[src/main/scala/chisel3/util/OneHot.scala 83:30]
  wire  _outSelRespVec_T = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _outSelRespVec_T_1 = state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 41:59]
  wire  _outSelRespVec_T_2 = _outSelRespVec_T & state == 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 41:50]
  reg  outSelRespVec_0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_2; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_3; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  reg  outSelRespVec_4; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire [4:0] _reqInvalidAddr_T = {outSelVec_4,outSelVec_3,outSelVec_2,outSelVec_1,outSelVec_0}; // @[src/main/scala/bus/simplebus/Crossbar.scala 42:54]
  wire  reqInvalidAddr = io_in_req_valid & ~(|_reqInvalidAddr_T); // @[src/main/scala/bus/simplebus/Crossbar.scala 42:40]
  wire  _T_7 = io_in_resp_ready & io_in_resp_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire [1:0] _GEN_7 = _T_7 ? 2'h0 : state; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22 56:{44,52}]
  wire  _io_in_req_ready_T_8 = outSelVec_0 & io_out_0_req_ready | outSelVec_1 & io_out_1_req_ready | outSelVec_2 &
    io_out_2_req_ready | outSelVec_3 & io_out_3_req_ready | outSelVec_4 & io_out_4_req_ready; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_in_resp_valid_T_8 = outSelRespVec_0 & io_out_0_resp_valid | outSelRespVec_1 & io_out_1_resp_valid |
    outSelRespVec_2 & io_out_2_resp_valid | outSelRespVec_3 & io_out_3_resp_valid | outSelRespVec_4 &
    io_out_4_resp_valid; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T = outSelRespVec_0 ? io_out_0_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_2 = outSelRespVec_2 ? io_out_2_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_3 = outSelRespVec_3 ? io_out_3_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_4 = outSelRespVec_4 ? io_out_4_resp_bits_rdata : 64'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_6 = _io_in_resp_bits_T | _io_in_resp_bits_T_2; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] _io_in_resp_bits_T_7 = _io_in_resp_bits_T_6 | _io_in_resp_bits_T_3; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_9 = outSelRespVec_0 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_10 = outSelRespVec_1 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_11 = outSelRespVec_2 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_12 = outSelRespVec_3 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_13 = outSelRespVec_4 ? 4'h6 : 4'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_14 = _io_in_resp_bits_T_9 | _io_in_resp_bits_T_10; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_15 = _io_in_resp_bits_T_14 | _io_in_resp_bits_T_11; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [3:0] _io_in_resp_bits_T_16 = _io_in_resp_bits_T_15 | _io_in_resp_bits_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [1:0] state_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
  wire [1:0] state_t = state ^ state_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
  wire  toggle_10811_clock;
  wire  toggle_10811_reset;
  wire [1:0] toggle_10811_valid;
  reg [1:0] toggle_10811_valid_reg;
  reg  outSelRespVec_0_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire  outSelRespVec_0_t = outSelRespVec_0 ^ outSelRespVec_0_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire  toggle_10813_clock;
  wire  toggle_10813_reset;
  wire  toggle_10813_valid;
  reg  toggle_10813_valid_reg;
  reg  outSelRespVec_1_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire  outSelRespVec_1_t = outSelRespVec_1 ^ outSelRespVec_1_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire  toggle_10814_clock;
  wire  toggle_10814_reset;
  wire  toggle_10814_valid;
  reg  toggle_10814_valid_reg;
  reg  outSelRespVec_2_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire  outSelRespVec_2_t = outSelRespVec_2 ^ outSelRespVec_2_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire  toggle_10815_clock;
  wire  toggle_10815_reset;
  wire  toggle_10815_valid;
  reg  toggle_10815_valid_reg;
  reg  outSelRespVec_3_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire  outSelRespVec_3_t = outSelRespVec_3 ^ outSelRespVec_3_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire  toggle_10816_clock;
  wire  toggle_10816_reset;
  wire  toggle_10816_valid;
  reg  toggle_10816_valid_reg;
  reg  outSelRespVec_4_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire  outSelRespVec_4_t = outSelRespVec_4 ^ outSelRespVec_4_p; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
  wire  toggle_10817_clock;
  wire  toggle_10817_reset;
  wire  toggle_10817_valid;
  reg  toggle_10817_valid_reg;
  GEN_w2_toggle #(.COVER_INDEX(10811)) toggle_10811 (
    .clock(toggle_10811_clock),
    .reset(toggle_10811_reset),
    .valid(toggle_10811_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10813)) toggle_10813 (
    .clock(toggle_10813_clock),
    .reset(toggle_10813_reset),
    .valid(toggle_10813_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10814)) toggle_10814 (
    .clock(toggle_10814_clock),
    .reset(toggle_10814_reset),
    .valid(toggle_10814_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10815)) toggle_10815 (
    .clock(toggle_10815_clock),
    .reset(toggle_10815_reset),
    .valid(toggle_10815_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10816)) toggle_10816 (
    .clock(toggle_10816_clock),
    .reset(toggle_10816_reset),
    .valid(toggle_10816_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10817)) toggle_10817 (
    .clock(toggle_10817_clock),
    .reset(toggle_10817_reset),
    .valid(toggle_10817_valid)
  );
  assign io_in_req_ready = _io_in_req_ready_T_8 | reqInvalidAddr; // @[src/main/scala/bus/simplebus/Crossbar.scala 61:64]
  assign io_in_resp_valid = _io_in_resp_valid_T_8 | state == 2'h2; // @[src/main/scala/bus/simplebus/Crossbar.scala 71:70]
  assign io_in_resp_bits_cmd = _io_in_resp_bits_T_16 | _io_in_resp_bits_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_in_resp_bits_rdata = _io_in_resp_bits_T_7 | _io_in_resp_bits_T_4; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  assign io_out_0_req_valid = outSelVec_0 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_0_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_0_resp_ready = outSelRespVec_0 & io_in_resp_ready & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_1_req_valid = outSelVec_1 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_1_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_1_resp_ready = outSelRespVec_1 & io_in_resp_ready & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_2_req_valid = outSelVec_2 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_2_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_2_resp_ready = outSelRespVec_2 & io_in_resp_ready & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_3_req_valid = outSelVec_3 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_3_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_3_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_3_resp_ready = outSelRespVec_3 & io_in_resp_ready & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign io_out_4_req_valid = outSelVec_4 & io_in_req_valid & _outSelRespVec_T_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 63:60]
  assign io_out_4_req_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_4_req_bits_cmd = io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_4_req_bits_wmask = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_4_req_bits_wdata = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/Crossbar.scala 64:24]
  assign io_out_4_resp_ready = outSelRespVec_4 & io_in_resp_ready & state == 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 69:66]
  assign toggle_10811_clock = clock;
  assign toggle_10811_reset = reset;
  assign toggle_10811_valid = state ^ toggle_10811_valid_reg;
  assign toggle_10813_clock = clock;
  assign toggle_10813_reset = reset;
  assign toggle_10813_valid = outSelRespVec_0 ^ toggle_10813_valid_reg;
  assign toggle_10814_clock = clock;
  assign toggle_10814_reset = reset;
  assign toggle_10814_valid = outSelRespVec_1 ^ toggle_10814_valid_reg;
  assign toggle_10815_clock = clock;
  assign toggle_10815_reset = reset;
  assign toggle_10815_valid = outSelRespVec_2 ^ toggle_10815_valid_reg;
  assign toggle_10816_clock = clock;
  assign toggle_10816_reset = reset;
  assign toggle_10816_valid = outSelRespVec_3 ^ toggle_10816_valid_reg;
  assign toggle_10817_clock = clock;
  assign toggle_10817_reset = reset;
  assign toggle_10817_valid = outSelRespVec_4 ^ toggle_10817_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
      state <= 2'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
    end else if (2'h0 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      if (reqInvalidAddr) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 54:29]
        state <= 2'h2; // @[src/main/scala/bus/simplebus/Crossbar.scala 54:37]
      end else if (_outSelRespVec_T) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 53:31]
        state <= 2'h1; // @[src/main/scala/bus/simplebus/Crossbar.scala 53:39]
      end
    end else if (2'h1 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      state <= _GEN_7;
    end else if (2'h2 == state) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 51:18]
      state <= _GEN_7;
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_0 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_0 <= outSelVec_0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_1 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_1 <= outSelVec_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_2 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_2 <= outSelVec_2; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_3 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_3 <= outSelVec_3; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    if (reset) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_4 <= 1'h0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end else if (_outSelRespVec_T_2) begin // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
      outSelRespVec_4 <= outSelVec_4; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~reqInvalidAddr)) begin
          $fwrite(32'h80000002,
            "Assertion failed: address decode error, bad addr = 0x%x\n\n    at Crossbar.scala:49 assert(!reqInvalidAddr, \"address decode error, bad addr = 0x%%%%x\\n\", addr)\n"
            ,io_in_req_bits_addr); // @[src/main/scala/bus/simplebus/Crossbar.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    state_p <= state; // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
    toggle_10811_valid_reg <= state;
    outSelRespVec_0_p <= outSelRespVec_0; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    toggle_10813_valid_reg <= outSelRespVec_0;
    outSelRespVec_1_p <= outSelRespVec_1; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    toggle_10814_valid_reg <= outSelRespVec_1;
    outSelRespVec_2_p <= outSelRespVec_2; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    toggle_10815_valid_reg <= outSelRespVec_2;
    outSelRespVec_3_p <= outSelRespVec_3; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    toggle_10816_valid_reg <= outSelRespVec_3;
    outSelRespVec_4_p <= outSelRespVec_4; // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    toggle_10817_valid_reg <= outSelRespVec_4;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  outSelRespVec_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  outSelRespVec_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  outSelRespVec_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  outSelRespVec_3 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  outSelRespVec_4 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  state_p = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  toggle_10811_valid_reg = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  outSelRespVec_0_p = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  toggle_10813_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  outSelRespVec_1_p = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  toggle_10814_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  outSelRespVec_2_p = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  toggle_10815_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  outSelRespVec_3_p = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  toggle_10816_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  outSelRespVec_4_p = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  toggle_10817_valid_reg = _RAND_17[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~reqInvalidAddr); // @[src/main/scala/bus/simplebus/Crossbar.scala 49:9]
    end
    //
    if (enToggle_past) begin
      cover(state_t[0]); // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(state_t[1]); // @[src/main/scala/bus/simplebus/Crossbar.scala 32:22]
    end
    //
    if (enToggle_past) begin
      cover(outSelRespVec_0_t); // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    //
    if (enToggle_past) begin
      cover(outSelRespVec_1_t); // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    //
    if (enToggle_past) begin
      cover(outSelRespVec_2_t); // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    //
    if (enToggle_past) begin
      cover(outSelRespVec_3_t); // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
    //
    if (enToggle_past) begin
      cover(outSelRespVec_4_t); // @[src/main/scala/bus/simplebus/Crossbar.scala 39:32]
    end
  end
endmodule
module AXI4UART(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_out_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [7:0]  io_extra_out_ch, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_in_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_extra_in_ch // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  wire  _r_busy_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _r_busy_T_1 = io_in_r_ready & io_in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _r_busy_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_2 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io_in_b_ready & io_in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _w_busy_T | _GEN_4; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [31:0] txfifo; // @[src/main/scala/device/AXI4UART.scala 29:19]
  reg [31:0] stat; // @[src/main/scala/device/AXI4UART.scala 30:21]
  reg [31:0] ctrl; // @[src/main/scala/device/AXI4UART.scala 31:21]
  wire  _io_extra_out_valid_T_1 = io_in_aw_bits_addr[3:0] == 4'h4; // @[src/main/scala/device/AXI4UART.scala 33:41]
  wire [7:0] _T_5 = io_in_w_bits_strb >> io_in_aw_bits_addr[2:0]; // @[src/main/scala/device/AXI4UART.scala 45:79]
  wire [7:0] _T_14 = _T_5[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_15 = _T_5[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_16 = _T_5[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_17 = _T_5[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_18 = _T_5[4] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_19 = _T_5[5] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_20 = _T_5[6] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_21 = _T_5[7] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [63:0] _T_22 = {_T_21,_T_20,_T_19,_T_18,_T_17,_T_16,_T_15,_T_14}; // @[src/main/scala/utils/BitUtils.scala 27:27]
  wire  _io_in_r_bits_data_T = 4'h0 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_1 = 4'h4 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_2 = 4'h8 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_3 = 4'hc == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [7:0] _io_in_r_bits_data_T_4 = _io_in_r_bits_data_T ? io_extra_in_ch : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_5 = _io_in_r_bits_data_T_1 ? txfifo : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_6 = _io_in_r_bits_data_T_2 ? stat : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_7 = _io_in_r_bits_data_T_3 ? ctrl : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _GEN_18 = {{24'd0}, _io_in_r_bits_data_T_4}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_8 = _GEN_18 | _io_in_r_bits_data_T_5; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_9 = _io_in_r_bits_data_T_8 | _io_in_r_bits_data_T_6; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_10 = _io_in_r_bits_data_T_9 | _io_in_r_bits_data_T_7; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _txfifo_T = io_in_w_bits_data[31:0] & _T_22[31:0]; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [31:0] _txfifo_T_1 = ~_T_22[31:0]; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [31:0] _txfifo_T_2 = txfifo & _txfifo_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _txfifo_T_3 = _txfifo_T | _txfifo_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _stat_T_2 = stat & _txfifo_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _stat_T_3 = _txfifo_T | _stat_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _ctrl_T_2 = ctrl & _txfifo_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _ctrl_T_3 = _txfifo_T | _ctrl_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  r_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  r_busy_t = r_busy ^ r_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10818_clock;
  wire  toggle_10818_reset;
  wire  toggle_10818_valid;
  reg  toggle_10818_valid_reg;
  reg  ren_REG_p; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  ren_REG_t = ren_REG ^ ren_REG_p; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  toggle_10819_clock;
  wire  toggle_10819_reset;
  wire  toggle_10819_valid;
  reg  toggle_10819_valid_reg;
  reg  io_in_r_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  io_in_r_valid_r_t = io_in_r_valid_r ^ io_in_r_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10820_clock;
  wire  toggle_10820_reset;
  wire  toggle_10820_valid;
  reg  toggle_10820_valid_reg;
  reg  w_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  w_busy_t = w_busy ^ w_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10821_clock;
  wire  toggle_10821_reset;
  wire  toggle_10821_valid;
  reg  toggle_10821_valid_reg;
  reg  io_in_b_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  io_in_b_valid_r_t = io_in_b_valid_r ^ io_in_b_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10822_clock;
  wire  toggle_10822_reset;
  wire  toggle_10822_valid;
  reg  toggle_10822_valid_reg;
  reg [31:0] txfifo_p; // @[src/main/scala/device/AXI4UART.scala 29:19]
  wire [31:0] txfifo_t = txfifo ^ txfifo_p; // @[src/main/scala/device/AXI4UART.scala 29:19]
  wire  toggle_10823_clock;
  wire  toggle_10823_reset;
  wire [31:0] toggle_10823_valid;
  reg [31:0] toggle_10823_valid_reg;
  reg [31:0] stat_p; // @[src/main/scala/device/AXI4UART.scala 30:21]
  wire [31:0] stat_t = stat ^ stat_p; // @[src/main/scala/device/AXI4UART.scala 30:21]
  wire  toggle_10855_clock;
  wire  toggle_10855_reset;
  wire [31:0] toggle_10855_valid;
  reg [31:0] toggle_10855_valid_reg;
  reg [31:0] ctrl_p; // @[src/main/scala/device/AXI4UART.scala 31:21]
  wire [31:0] ctrl_t = ctrl ^ ctrl_p; // @[src/main/scala/device/AXI4UART.scala 31:21]
  wire  toggle_10887_clock;
  wire  toggle_10887_reset;
  wire [31:0] toggle_10887_valid;
  reg [31:0] toggle_10887_valid_reg;
  GEN_w1_toggle #(.COVER_INDEX(10818)) toggle_10818 (
    .clock(toggle_10818_clock),
    .reset(toggle_10818_reset),
    .valid(toggle_10818_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10819)) toggle_10819 (
    .clock(toggle_10819_clock),
    .reset(toggle_10819_reset),
    .valid(toggle_10819_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10820)) toggle_10820 (
    .clock(toggle_10820_clock),
    .reset(toggle_10820_reset),
    .valid(toggle_10820_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10821)) toggle_10821 (
    .clock(toggle_10821_clock),
    .reset(toggle_10821_reset),
    .valid(toggle_10821_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10822)) toggle_10822 (
    .clock(toggle_10822_clock),
    .reset(toggle_10822_reset),
    .valid(toggle_10822_valid)
  );
  GEN_w32_toggle #(.COVER_INDEX(10823)) toggle_10823 (
    .clock(toggle_10823_clock),
    .reset(toggle_10823_reset),
    .valid(toggle_10823_valid)
  );
  GEN_w32_toggle #(.COVER_INDEX(10855)) toggle_10855 (
    .clock(toggle_10855_clock),
    .reset(toggle_10855_reset),
    .valid(toggle_10855_valid)
  );
  GEN_w32_toggle #(.COVER_INDEX(10887)) toggle_10887 (
    .clock(toggle_10887_clock),
    .reset(toggle_10887_reset),
    .valid(toggle_10887_valid)
  );
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = {{32'd0}, _io_in_r_bits_data_T_10}; // @[src/main/scala/utils/RegMap.scala 30:11]
  assign io_extra_out_valid = io_in_aw_bits_addr[3:0] == 4'h4 & _io_in_b_valid_T; // @[src/main/scala/device/AXI4UART.scala 33:49]
  assign io_extra_out_ch = io_in_w_bits_data[7:0]; // @[src/main/scala/device/AXI4UART.scala 34:40]
  assign io_extra_in_valid = io_in_ar_bits_addr[3:0] == 4'h0 & _r_busy_T_1; // @[src/main/scala/device/AXI4UART.scala 35:48]
  assign toggle_10818_clock = clock;
  assign toggle_10818_reset = reset;
  assign toggle_10818_valid = r_busy ^ toggle_10818_valid_reg;
  assign toggle_10819_clock = clock;
  assign toggle_10819_reset = reset;
  assign toggle_10819_valid = ren_REG ^ toggle_10819_valid_reg;
  assign toggle_10820_clock = clock;
  assign toggle_10820_reset = reset;
  assign toggle_10820_valid = io_in_r_valid_r ^ toggle_10820_valid_reg;
  assign toggle_10821_clock = clock;
  assign toggle_10821_reset = reset;
  assign toggle_10821_valid = w_busy ^ toggle_10821_valid_reg;
  assign toggle_10822_clock = clock;
  assign toggle_10822_reset = reset;
  assign toggle_10822_valid = io_in_b_valid_r ^ toggle_10822_valid_reg;
  assign toggle_10823_clock = clock;
  assign toggle_10823_reset = reset;
  assign toggle_10823_valid = txfifo ^ toggle_10823_valid_reg;
  assign toggle_10855_clock = clock;
  assign toggle_10855_reset = reset;
  assign toggle_10855_valid = stat ^ toggle_10855_valid_reg;
  assign toggle_10887_clock = clock;
  assign toggle_10887_reset = reset;
  assign toggle_10887_valid = ctrl ^ toggle_10887_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
    if (_io_in_b_valid_T & _io_extra_out_valid_T_1) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      txfifo <= _txfifo_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4UART.scala 30:21]
      stat <= 32'h1; // @[src/main/scala/device/AXI4UART.scala 30:21]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[3:0] == 4'h8) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      stat <= _stat_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4UART.scala 31:21]
      ctrl <= 32'h0; // @[src/main/scala/device/AXI4UART.scala 31:21]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[3:0] == 4'hc) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      ctrl <= _ctrl_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    r_busy_p <= r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10818_valid_reg <= r_busy;
    ren_REG_p <= ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    toggle_10819_valid_reg <= ren_REG;
    io_in_r_valid_r_p <= io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10820_valid_reg <= io_in_r_valid_r;
    w_busy_p <= w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10821_valid_reg <= w_busy;
    io_in_b_valid_r_p <= io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10822_valid_reg <= io_in_b_valid_r;
    txfifo_p <= txfifo; // @[src/main/scala/device/AXI4UART.scala 29:19]
    toggle_10823_valid_reg <= txfifo;
    stat_p <= stat; // @[src/main/scala/device/AXI4UART.scala 30:21]
    toggle_10855_valid_reg <= stat;
    ctrl_p <= ctrl; // @[src/main/scala/device/AXI4UART.scala 31:21]
    toggle_10887_valid_reg <= ctrl;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  txfifo = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  stat = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  ctrl = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  r_busy_p = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  toggle_10818_valid_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ren_REG_p = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  toggle_10819_valid_reg = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  io_in_r_valid_r_p = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  toggle_10820_valid_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  w_busy_p = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  toggle_10821_valid_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  io_in_b_valid_r_p = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  toggle_10822_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  txfifo_p = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  toggle_10823_valid_reg = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  stat_p = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  toggle_10855_valid_reg = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  ctrl_p = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  toggle_10887_valid_reg = _RAND_23[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(r_busy_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(ren_REG_t); // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_valid_r_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(w_busy_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(io_in_b_valid_r_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[0]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[1]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[2]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[3]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[4]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[5]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[6]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[7]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[8]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[9]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[10]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[11]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[12]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[13]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[14]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[15]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[16]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[17]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[18]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[19]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[20]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[21]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[22]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[23]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[24]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[25]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[26]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[27]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[28]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[29]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[30]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(txfifo_t[31]); // @[src/main/scala/device/AXI4UART.scala 29:19]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[0]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[1]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[2]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[3]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[4]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[5]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[6]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[7]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[8]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[9]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[10]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[11]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[12]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[13]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[14]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[15]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[16]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[17]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[18]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[19]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[20]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[21]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[22]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[23]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[24]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[25]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[26]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[27]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[28]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[29]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[30]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(stat_t[31]); // @[src/main/scala/device/AXI4UART.scala 30:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[0]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[1]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[2]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[3]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[4]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[5]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[6]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[7]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[8]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[9]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[10]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[11]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[12]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[13]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[14]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[15]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[16]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[17]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[18]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[19]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[20]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[21]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[22]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[23]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[24]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[25]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[26]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[27]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[28]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[29]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[30]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
    //
    if (enToggle_past) begin
      cover(ctrl_t[31]); // @[src/main/scala/device/AXI4UART.scala 31:21]
    end
  end
endmodule
module VGACtrl(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_extra_sync // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire  _r_busy_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _r_busy_T_1 = io_in_r_ready & io_in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _r_busy_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_2 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io_in_b_ready & io_in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _w_busy_T | _GEN_4; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_r_bits_data_T = 4'h0 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _io_in_r_bits_data_T_1 = 4'h4 == io_in_ar_bits_addr[3:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _io_in_r_bits_data_T_2 = _io_in_r_bits_data_T ? 32'h190012c : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire  _io_in_r_bits_data_T_3 = _io_in_r_bits_data_T_1 & _w_busy_T; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _GEN_13 = {{31'd0}, _io_in_r_bits_data_T_3}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _io_in_r_bits_data_T_4 = _io_in_r_bits_data_T_2 | _GEN_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  r_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  r_busy_t = r_busy ^ r_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10919_clock;
  wire  toggle_10919_reset;
  wire  toggle_10919_valid;
  reg  toggle_10919_valid_reg;
  reg  ren_REG_p; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  ren_REG_t = ren_REG ^ ren_REG_p; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  toggle_10920_clock;
  wire  toggle_10920_reset;
  wire  toggle_10920_valid;
  reg  toggle_10920_valid_reg;
  reg  io_in_r_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  io_in_r_valid_r_t = io_in_r_valid_r ^ io_in_r_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10921_clock;
  wire  toggle_10921_reset;
  wire  toggle_10921_valid;
  reg  toggle_10921_valid_reg;
  reg  w_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  w_busy_t = w_busy ^ w_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10922_clock;
  wire  toggle_10922_reset;
  wire  toggle_10922_valid;
  reg  toggle_10922_valid_reg;
  reg  io_in_b_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  io_in_b_valid_r_t = io_in_b_valid_r ^ io_in_b_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10923_clock;
  wire  toggle_10923_reset;
  wire  toggle_10923_valid;
  reg  toggle_10923_valid_reg;
  GEN_w1_toggle #(.COVER_INDEX(10919)) toggle_10919 (
    .clock(toggle_10919_clock),
    .reset(toggle_10919_reset),
    .valid(toggle_10919_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10920)) toggle_10920 (
    .clock(toggle_10920_clock),
    .reset(toggle_10920_reset),
    .valid(toggle_10920_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10921)) toggle_10921 (
    .clock(toggle_10921_clock),
    .reset(toggle_10921_reset),
    .valid(toggle_10921_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10922)) toggle_10922 (
    .clock(toggle_10922_clock),
    .reset(toggle_10922_reset),
    .valid(toggle_10922_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10923)) toggle_10923 (
    .clock(toggle_10923_clock),
    .reset(toggle_10923_reset),
    .valid(toggle_10923_valid)
  );
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = {{32'd0}, _io_in_r_bits_data_T_4}; // @[src/main/scala/utils/RegMap.scala 30:11]
  assign io_extra_sync = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  assign toggle_10919_clock = clock;
  assign toggle_10919_reset = reset;
  assign toggle_10919_valid = r_busy ^ toggle_10919_valid_reg;
  assign toggle_10920_clock = clock;
  assign toggle_10920_reset = reset;
  assign toggle_10920_valid = ren_REG ^ toggle_10920_valid_reg;
  assign toggle_10921_clock = clock;
  assign toggle_10921_reset = reset;
  assign toggle_10921_valid = io_in_r_valid_r ^ toggle_10921_valid_reg;
  assign toggle_10922_clock = clock;
  assign toggle_10922_reset = reset;
  assign toggle_10922_valid = w_busy ^ toggle_10922_valid_reg;
  assign toggle_10923_clock = clock;
  assign toggle_10923_reset = reset;
  assign toggle_10923_valid = io_in_b_valid_r ^ toggle_10923_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    r_busy_p <= r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10919_valid_reg <= r_busy;
    ren_REG_p <= ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    toggle_10920_valid_reg <= ren_REG;
    io_in_r_valid_r_p <= io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10921_valid_reg <= io_in_r_valid_r;
    w_busy_p <= w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10922_valid_reg <= w_busy;
    io_in_b_valid_r_p <= io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10923_valid_reg <= io_in_b_valid_r;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  r_busy_p = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  toggle_10919_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  ren_REG_p = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  toggle_10920_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  io_in_r_valid_r_p = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  toggle_10921_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  w_busy_p = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  toggle_10922_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  io_in_b_valid_r_p = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  toggle_10923_valid_reg = _RAND_14[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(r_busy_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(ren_REG_t); // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_valid_r_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(w_busy_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(io_in_b_valid_r_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
  end
endmodule
module AXI4RAM_1(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] rdata_mem_0 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_0_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_0_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_0_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_0_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_0_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_0_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_0_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_1 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_1_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_1_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_1_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_1_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_1_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_1_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_1_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_2 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_2_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_2_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_2_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_2_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_2_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_2_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_2_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_3 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_3_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_3_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_3_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_3_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_3_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_3_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_3_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_4 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_4_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_4_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_4_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_4_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_4_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_4_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_4_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_5 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_5_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_5_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_5_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_5_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_5_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_5_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_5_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_6 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_6_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_6_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_6_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_6_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_6_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_6_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_6_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  reg [7:0] rdata_mem_7 [0:59999]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_7_rdata_MPORT_1_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_7_rdata_MPORT_1_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_7_rdata_MPORT_1_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [7:0] rdata_mem_7_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire [15:0] rdata_mem_7_rdata_MPORT_addr; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_7_rdata_MPORT_mask; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  rdata_mem_7_rdata_MPORT_en; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  wire  _r_busy_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = io_in_r_valid ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _r_busy_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_2 = io_in_r_valid ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io_in_b_ready & io_in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _w_busy_T | _GEN_4; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire [31:0] _wIdx_T = io_in_aw_bits_addr & 32'h7ffff; // @[src/main/scala/device/AXI4RAM.scala 32:33]
  wire [29:0] _wIdx_T_2 = {{1'd0}, _wIdx_T[31:3]}; // @[src/main/scala/device/AXI4RAM.scala 35:27]
  wire [28:0] wIdx = _wIdx_T_2[28:0]; // @[src/main/scala/device/AXI4RAM.scala 35:27]
  wire [31:0] _rIdx_T = io_in_ar_bits_addr & 32'h7ffff; // @[src/main/scala/device/AXI4RAM.scala 32:33]
  wire [29:0] _rIdx_T_2 = {{1'd0}, _rIdx_T[31:3]}; // @[src/main/scala/device/AXI4RAM.scala 36:27]
  wire [28:0] rIdx = _rIdx_T_2[28:0]; // @[src/main/scala/device/AXI4RAM.scala 36:27]
  wire  _wen_T_1 = wIdx < 29'hea60; // @[src/main/scala/device/AXI4RAM.scala 33:32]
  wire [63:0] _rdata_T_12 = {rdata_mem_7_rdata_MPORT_1_data,rdata_mem_6_rdata_MPORT_1_data,
    rdata_mem_5_rdata_MPORT_1_data,rdata_mem_4_rdata_MPORT_1_data,rdata_mem_3_rdata_MPORT_1_data,
    rdata_mem_2_rdata_MPORT_1_data,rdata_mem_1_rdata_MPORT_1_data,rdata_mem_0_rdata_MPORT_1_data}; // @[src/main/scala/device/AXI4RAM.scala 55:18]
  reg [63:0] rdata; // @[src/main/scala/device/AXI4RAM.scala 55:14]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  r_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  r_busy_t = r_busy ^ r_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10924_clock;
  wire  toggle_10924_reset;
  wire  toggle_10924_valid;
  reg  toggle_10924_valid_reg;
  reg  ren_REG_p; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  ren_REG_t = ren_REG ^ ren_REG_p; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  toggle_10925_clock;
  wire  toggle_10925_reset;
  wire  toggle_10925_valid;
  reg  toggle_10925_valid_reg;
  reg  io_in_r_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  io_in_r_valid_r_t = io_in_r_valid_r ^ io_in_r_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10926_clock;
  wire  toggle_10926_reset;
  wire  toggle_10926_valid;
  reg  toggle_10926_valid_reg;
  reg  w_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  w_busy_t = w_busy ^ w_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10927_clock;
  wire  toggle_10927_reset;
  wire  toggle_10927_valid;
  reg  toggle_10927_valid_reg;
  reg  io_in_b_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  io_in_b_valid_r_t = io_in_b_valid_r ^ io_in_b_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10928_clock;
  wire  toggle_10928_reset;
  wire  toggle_10928_valid;
  reg  toggle_10928_valid_reg;
  reg [63:0] rdata_p; // @[src/main/scala/device/AXI4RAM.scala 55:14]
  wire [63:0] rdata_t = rdata ^ rdata_p; // @[src/main/scala/device/AXI4RAM.scala 55:14]
  wire  toggle_10929_clock;
  wire  toggle_10929_reset;
  wire [63:0] toggle_10929_valid;
  reg [63:0] toggle_10929_valid_reg;
  GEN_w1_toggle #(.COVER_INDEX(10924)) toggle_10924 (
    .clock(toggle_10924_clock),
    .reset(toggle_10924_reset),
    .valid(toggle_10924_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10925)) toggle_10925 (
    .clock(toggle_10925_clock),
    .reset(toggle_10925_reset),
    .valid(toggle_10925_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10926)) toggle_10926 (
    .clock(toggle_10926_clock),
    .reset(toggle_10926_reset),
    .valid(toggle_10926_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10927)) toggle_10927 (
    .clock(toggle_10927_clock),
    .reset(toggle_10927_reset),
    .valid(toggle_10927_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(10928)) toggle_10928 (
    .clock(toggle_10928_clock),
    .reset(toggle_10928_reset),
    .valid(toggle_10928_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(10929)) toggle_10929 (
    .clock(toggle_10929_clock),
    .reset(toggle_10929_reset),
    .valid(toggle_10929_valid)
  );
  assign rdata_mem_0_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_0_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_0_rdata_MPORT_1_data = rdata_mem_0[rdata_mem_0_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_0_rdata_MPORT_1_data = rdata_mem_0_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_1[7:0] :
    rdata_mem_0[rdata_mem_0_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_0_rdata_MPORT_data = io_in_w_bits_data[7:0];
  assign rdata_mem_0_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_0_rdata_MPORT_mask = io_in_w_bits_strb[0];
  assign rdata_mem_0_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_1_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_1_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_1_rdata_MPORT_1_data = rdata_mem_1[rdata_mem_1_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_1_rdata_MPORT_1_data = rdata_mem_1_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_3[7:0] :
    rdata_mem_1[rdata_mem_1_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_1_rdata_MPORT_data = io_in_w_bits_data[15:8];
  assign rdata_mem_1_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_1_rdata_MPORT_mask = io_in_w_bits_strb[1];
  assign rdata_mem_1_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_2_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_2_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_2_rdata_MPORT_1_data = rdata_mem_2[rdata_mem_2_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_2_rdata_MPORT_1_data = rdata_mem_2_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_5[7:0] :
    rdata_mem_2[rdata_mem_2_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_2_rdata_MPORT_data = io_in_w_bits_data[23:16];
  assign rdata_mem_2_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_2_rdata_MPORT_mask = io_in_w_bits_strb[2];
  assign rdata_mem_2_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_3_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_3_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_3_rdata_MPORT_1_data = rdata_mem_3[rdata_mem_3_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_3_rdata_MPORT_1_data = rdata_mem_3_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_7[7:0] :
    rdata_mem_3[rdata_mem_3_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_3_rdata_MPORT_data = io_in_w_bits_data[31:24];
  assign rdata_mem_3_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_3_rdata_MPORT_mask = io_in_w_bits_strb[3];
  assign rdata_mem_3_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_4_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_4_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_4_rdata_MPORT_1_data = rdata_mem_4[rdata_mem_4_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_4_rdata_MPORT_1_data = rdata_mem_4_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_9[7:0] :
    rdata_mem_4[rdata_mem_4_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_4_rdata_MPORT_data = io_in_w_bits_data[39:32];
  assign rdata_mem_4_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_4_rdata_MPORT_mask = io_in_w_bits_strb[4];
  assign rdata_mem_4_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_5_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_5_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_5_rdata_MPORT_1_data = rdata_mem_5[rdata_mem_5_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_5_rdata_MPORT_1_data = rdata_mem_5_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_11[7:0] :
    rdata_mem_5[rdata_mem_5_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_5_rdata_MPORT_data = io_in_w_bits_data[47:40];
  assign rdata_mem_5_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_5_rdata_MPORT_mask = io_in_w_bits_strb[5];
  assign rdata_mem_5_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_6_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_6_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_6_rdata_MPORT_1_data = rdata_mem_6[rdata_mem_6_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_6_rdata_MPORT_1_data = rdata_mem_6_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_13[7:0] :
    rdata_mem_6[rdata_mem_6_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_6_rdata_MPORT_data = io_in_w_bits_data[55:48];
  assign rdata_mem_6_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_6_rdata_MPORT_mask = io_in_w_bits_strb[6];
  assign rdata_mem_6_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign rdata_mem_7_rdata_MPORT_1_en = 1'h1;
  assign rdata_mem_7_rdata_MPORT_1_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_7_rdata_MPORT_1_data = rdata_mem_7[rdata_mem_7_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `else
  assign rdata_mem_7_rdata_MPORT_1_data = rdata_mem_7_rdata_MPORT_1_addr >= 16'hea60 ? _RAND_15[7:0] :
    rdata_mem_7[rdata_mem_7_rdata_MPORT_1_addr]; // @[src/main/scala/device/AXI4RAM.scala 50:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rdata_mem_7_rdata_MPORT_data = io_in_w_bits_data[63:56];
  assign rdata_mem_7_rdata_MPORT_addr = wIdx[15:0];
  assign rdata_mem_7_rdata_MPORT_mask = io_in_w_bits_strb[7];
  assign rdata_mem_7_rdata_MPORT_en = _io_in_b_valid_T & _wen_T_1;
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = 1'h1; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = rdata; // @[src/main/scala/device/AXI4RAM.scala 58:18]
  assign toggle_10924_clock = clock;
  assign toggle_10924_reset = reset;
  assign toggle_10924_valid = r_busy ^ toggle_10924_valid_reg;
  assign toggle_10925_clock = clock;
  assign toggle_10925_reset = reset;
  assign toggle_10925_valid = ren_REG ^ toggle_10925_valid_reg;
  assign toggle_10926_clock = clock;
  assign toggle_10926_reset = reset;
  assign toggle_10926_valid = io_in_r_valid_r ^ toggle_10926_valid_reg;
  assign toggle_10927_clock = clock;
  assign toggle_10927_reset = reset;
  assign toggle_10927_valid = w_busy ^ toggle_10927_valid_reg;
  assign toggle_10928_clock = clock;
  assign toggle_10928_reset = reset;
  assign toggle_10928_valid = io_in_b_valid_r ^ toggle_10928_valid_reg;
  assign toggle_10929_clock = clock;
  assign toggle_10929_reset = reset;
  assign toggle_10929_valid = rdata ^ toggle_10929_valid_reg;
  always @(posedge clock) begin
    if (rdata_mem_0_rdata_MPORT_en & rdata_mem_0_rdata_MPORT_mask) begin
      rdata_mem_0[rdata_mem_0_rdata_MPORT_addr] <= rdata_mem_0_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_1_rdata_MPORT_en & rdata_mem_1_rdata_MPORT_mask) begin
      rdata_mem_1[rdata_mem_1_rdata_MPORT_addr] <= rdata_mem_1_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_2_rdata_MPORT_en & rdata_mem_2_rdata_MPORT_mask) begin
      rdata_mem_2[rdata_mem_2_rdata_MPORT_addr] <= rdata_mem_2_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_3_rdata_MPORT_en & rdata_mem_3_rdata_MPORT_mask) begin
      rdata_mem_3[rdata_mem_3_rdata_MPORT_addr] <= rdata_mem_3_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_4_rdata_MPORT_en & rdata_mem_4_rdata_MPORT_mask) begin
      rdata_mem_4[rdata_mem_4_rdata_MPORT_addr] <= rdata_mem_4_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_5_rdata_MPORT_en & rdata_mem_5_rdata_MPORT_mask) begin
      rdata_mem_5[rdata_mem_5_rdata_MPORT_addr] <= rdata_mem_5_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_6_rdata_MPORT_en & rdata_mem_6_rdata_MPORT_mask) begin
      rdata_mem_6[rdata_mem_6_rdata_MPORT_addr] <= rdata_mem_6_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (rdata_mem_7_rdata_MPORT_en & rdata_mem_7_rdata_MPORT_mask) begin
      rdata_mem_7[rdata_mem_7_rdata_MPORT_addr] <= rdata_mem_7_rdata_MPORT_data; // @[src/main/scala/device/AXI4RAM.scala 50:18]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
    if (ren_REG) begin // @[src/main/scala/device/AXI4RAM.scala 55:14]
      rdata <= _rdata_T_12; // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    r_busy_p <= r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10924_valid_reg <= r_busy;
    ren_REG_p <= ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    toggle_10925_valid_reg <= ren_REG;
    io_in_r_valid_r_p <= io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10926_valid_reg <= io_in_r_valid_r;
    w_busy_p <= w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10927_valid_reg <= w_busy;
    io_in_b_valid_r_p <= io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10928_valid_reg <= io_in_b_valid_r;
    rdata_p <= rdata; // @[src/main/scala/device/AXI4RAM.scala 55:14]
    toggle_10929_valid_reg <= rdata;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {1{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
  _RAND_9 = {1{`RANDOM}};
  _RAND_11 = {1{`RANDOM}};
  _RAND_13 = {1{`RANDOM}};
  _RAND_15 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_0[initvar] = _RAND_0[7:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_1[initvar] = _RAND_2[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_2[initvar] = _RAND_4[7:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_3[initvar] = _RAND_6[7:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_4[initvar] = _RAND_8[7:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_5[initvar] = _RAND_10[7:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_6[initvar] = _RAND_12[7:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    rdata_mem_7[initvar] = _RAND_14[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  r_busy = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  ren_REG = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  w_busy = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  rdata = _RAND_21[63:0];
  _RAND_22 = {1{`RANDOM}};
  r_busy_p = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  toggle_10924_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  ren_REG_p = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  toggle_10925_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  io_in_r_valid_r_p = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  toggle_10926_valid_reg = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  w_busy_p = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  toggle_10927_valid_reg = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  io_in_b_valid_r_p = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  toggle_10928_valid_reg = _RAND_31[0:0];
  _RAND_32 = {2{`RANDOM}};
  rdata_p = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  toggle_10929_valid_reg = _RAND_33[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(r_busy_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(ren_REG_t); // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_valid_r_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(w_busy_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(io_in_b_valid_r_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[0]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[1]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[2]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[3]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[4]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[5]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[6]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[7]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[8]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[9]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[10]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[11]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[12]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[13]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[14]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[15]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[16]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[17]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[18]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[19]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[20]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[21]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[22]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[23]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[24]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[25]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[26]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[27]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[28]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[29]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[30]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[31]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[32]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[33]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[34]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[35]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[36]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[37]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[38]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[39]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[40]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[41]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[42]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[43]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[44]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[45]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[46]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[47]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[48]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[49]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[50]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[51]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[52]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[53]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[54]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[55]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[56]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[57]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[58]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[59]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[60]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[61]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[62]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
    //
    if (enToggle_past) begin
      cover(rdata_t[63]); // @[src/main/scala/device/AXI4RAM.scala 55:14]
    end
  end
endmodule
module AXI4VGA(
  input         clock,
  input         reset,
  output        io_in_fb_aw_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_fb_aw_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input  [31:0] io_in_fb_aw_bits_addr, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_fb_w_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_fb_w_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input  [63:0] io_in_fb_w_bits_data, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input  [7:0]  io_in_fb_w_bits_strb, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_fb_b_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_fb_b_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_fb_ar_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_fb_ar_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_fb_r_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_fb_r_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_ctrl_aw_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_ctrl_aw_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_ctrl_w_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_ctrl_w_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_ctrl_b_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_ctrl_b_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_ctrl_ar_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_ctrl_ar_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input  [31:0] io_in_ctrl_ar_bits_addr, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  input         io_in_ctrl_r_ready, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_in_ctrl_r_valid, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output [63:0] io_in_ctrl_r_bits_data, // @[src/main/scala/device/AXI4VGA.scala 117:14]
  output        io_vga_valid // @[src/main/scala/device/AXI4VGA.scala 117:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire  ctrl_clock; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_reset; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_aw_ready; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_aw_valid; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_w_ready; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_w_valid; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_b_ready; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_b_valid; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_ar_ready; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_ar_valid; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire [31:0] ctrl_io_in_ar_bits_addr; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_r_ready; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_in_r_valid; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire [63:0] ctrl_io_in_r_bits_data; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  ctrl_io_extra_sync; // @[src/main/scala/device/AXI4VGA.scala 125:20]
  wire  fb_clock; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_reset; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_aw_ready; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_aw_valid; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire [31:0] fb_io_in_aw_bits_addr; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_w_ready; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_w_valid; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire [63:0] fb_io_in_w_bits_data; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire [7:0] fb_io_in_w_bits_strb; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_b_ready; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_b_valid; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_ar_ready; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_ar_valid; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire [31:0] fb_io_in_ar_bits_addr; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_r_ready; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fb_io_in_r_valid; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire [63:0] fb_io_in_r_bits_data; // @[src/main/scala/device/AXI4VGA.scala 127:18]
  wire  fbHelper_clk; // @[src/main/scala/device/AXI4VGA.scala 171:26]
  wire  fbHelper_valid; // @[src/main/scala/device/AXI4VGA.scala 171:26]
  wire [31:0] fbHelper_pixel; // @[src/main/scala/device/AXI4VGA.scala 171:26]
  wire  fbHelper_sync; // @[src/main/scala/device/AXI4VGA.scala 171:26]
  wire  _io_in_fb_r_valid_T = io_in_fb_ar_ready & io_in_fb_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _io_in_fb_r_valid_T_1 = io_in_fb_r_ready & io_in_fb_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_fb_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _io_in_fb_r_valid_T_1 ? 1'h0 : io_in_fb_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _io_in_fb_r_valid_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [10:0] hCounter; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  wrap_wrap = hCounter == 11'h41f; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [10:0] _wrap_value_T_1 = hCounter + 11'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  reg [9:0] vCounter; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  wrap_wrap_1 = vCounter == 10'h273; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [9:0] _wrap_value_T_3 = vCounter + 10'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  hInRange = hCounter >= 11'ha8 & hCounter < 11'h3c8; // @[src/main/scala/device/AXI4VGA.scala 138:63]
  wire  vInRange = vCounter >= 10'h5 & vCounter < 10'h25d; // @[src/main/scala/device/AXI4VGA.scala 138:63]
  wire  hCounterIsOdd = hCounter[0]; // @[src/main/scala/device/AXI4VGA.scala 150:31]
  wire  hCounterIs2 = hCounter[1:0] == 2'h2; // @[src/main/scala/device/AXI4VGA.scala 151:35]
  wire  vCounterIsOdd = vCounter[0]; // @[src/main/scala/device/AXI4VGA.scala 152:31]
  wire  _nextPixel_T_2 = hCounter >= 11'ha7 & hCounter < 11'h3c7; // @[src/main/scala/device/AXI4VGA.scala 138:63]
  wire  nextPixel = _nextPixel_T_2 & vInRange & hCounterIsOdd; // @[src/main/scala/device/AXI4VGA.scala 155:78]
  wire  _fbPixelAddrV0_T_1 = nextPixel & ~vCounterIsOdd; // @[src/main/scala/device/AXI4VGA.scala 156:41]
  reg [16:0] fbPixelAddrV0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  fbPixelAddrV0_wrap_wrap = fbPixelAddrV0 == 17'h1d4bf; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [16:0] _fbPixelAddrV0_wrap_value_T_1 = fbPixelAddrV0 + 17'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire  _fbPixelAddrV1_T = nextPixel & vCounterIsOdd; // @[src/main/scala/device/AXI4VGA.scala 157:41]
  reg [16:0] fbPixelAddrV1; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  fbPixelAddrV1_wrap_wrap = fbPixelAddrV1 == 17'h1d4bf; // @[src/main/scala/chisel3/util/Counter.scala 73:24]
  wire [16:0] _fbPixelAddrV1_wrap_value_T_1 = fbPixelAddrV1 + 17'h1; // @[src/main/scala/chisel3/util/Counter.scala 77:24]
  wire [16:0] _fb_io_in_ar_bits_addr_T = vCounterIsOdd ? fbPixelAddrV1 : fbPixelAddrV0; // @[src/main/scala/device/AXI4VGA.scala 161:35]
  wire [18:0] _fb_io_in_ar_bits_addr_T_1 = {_fb_io_in_ar_bits_addr_T,2'h0}; // @[src/main/scala/device/AXI4VGA.scala 161:31]
  reg  fb_io_in_ar_valid_REG; // @[src/main/scala/device/AXI4VGA.scala 162:31]
  wire  _data_T = fb_io_in_r_ready & fb_io_in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg [63:0] data_r; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [63:0] _GEN_14 = _data_T ? fb_io_in_r_bits_data : data_r; // @[src/main/scala/utils/Hold.scala 23:{65,65,65}]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  io_in_fb_r_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  io_in_fb_r_valid_r_t = io_in_fb_r_valid_r ^ io_in_fb_r_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_10993_clock;
  wire  toggle_10993_reset;
  wire  toggle_10993_valid;
  reg  toggle_10993_valid_reg;
  reg [10:0] hCounter_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [10:0] hCounter_t = hCounter ^ hCounter_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  toggle_10994_clock;
  wire  toggle_10994_reset;
  wire [10:0] toggle_10994_valid;
  reg [10:0] toggle_10994_valid_reg;
  reg [9:0] vCounter_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [9:0] vCounter_t = vCounter ^ vCounter_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  toggle_11005_clock;
  wire  toggle_11005_reset;
  wire [9:0] toggle_11005_valid;
  reg [9:0] toggle_11005_valid_reg;
  reg [16:0] fbPixelAddrV0_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [16:0] fbPixelAddrV0_t = fbPixelAddrV0 ^ fbPixelAddrV0_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  toggle_11015_clock;
  wire  toggle_11015_reset;
  wire [16:0] toggle_11015_valid;
  reg [16:0] toggle_11015_valid_reg;
  reg [16:0] fbPixelAddrV1_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire [16:0] fbPixelAddrV1_t = fbPixelAddrV1 ^ fbPixelAddrV1_p; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
  wire  toggle_11032_clock;
  wire  toggle_11032_reset;
  wire [16:0] toggle_11032_valid;
  reg [16:0] toggle_11032_valid_reg;
  reg  fb_io_in_ar_valid_REG_p; // @[src/main/scala/device/AXI4VGA.scala 162:31]
  wire  fb_io_in_ar_valid_REG_t = fb_io_in_ar_valid_REG ^ fb_io_in_ar_valid_REG_p; // @[src/main/scala/device/AXI4VGA.scala 162:31]
  wire  toggle_11049_clock;
  wire  toggle_11049_reset;
  wire  toggle_11049_valid;
  reg  toggle_11049_valid_reg;
  reg [63:0] data_r_p; // @[src/main/scala/utils/Hold.scala 23:65]
  wire [63:0] data_r_t = data_r ^ data_r_p; // @[src/main/scala/utils/Hold.scala 23:65]
  wire  toggle_11050_clock;
  wire  toggle_11050_reset;
  wire [63:0] toggle_11050_valid;
  reg [63:0] toggle_11050_valid_reg;
  VGACtrl ctrl ( // @[src/main/scala/device/AXI4VGA.scala 125:20]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_in_aw_ready(ctrl_io_in_aw_ready),
    .io_in_aw_valid(ctrl_io_in_aw_valid),
    .io_in_w_ready(ctrl_io_in_w_ready),
    .io_in_w_valid(ctrl_io_in_w_valid),
    .io_in_b_ready(ctrl_io_in_b_ready),
    .io_in_b_valid(ctrl_io_in_b_valid),
    .io_in_ar_ready(ctrl_io_in_ar_ready),
    .io_in_ar_valid(ctrl_io_in_ar_valid),
    .io_in_ar_bits_addr(ctrl_io_in_ar_bits_addr),
    .io_in_r_ready(ctrl_io_in_r_ready),
    .io_in_r_valid(ctrl_io_in_r_valid),
    .io_in_r_bits_data(ctrl_io_in_r_bits_data),
    .io_extra_sync(ctrl_io_extra_sync)
  );
  AXI4RAM_1 fb ( // @[src/main/scala/device/AXI4VGA.scala 127:18]
    .clock(fb_clock),
    .reset(fb_reset),
    .io_in_aw_ready(fb_io_in_aw_ready),
    .io_in_aw_valid(fb_io_in_aw_valid),
    .io_in_aw_bits_addr(fb_io_in_aw_bits_addr),
    .io_in_w_ready(fb_io_in_w_ready),
    .io_in_w_valid(fb_io_in_w_valid),
    .io_in_w_bits_data(fb_io_in_w_bits_data),
    .io_in_w_bits_strb(fb_io_in_w_bits_strb),
    .io_in_b_ready(fb_io_in_b_ready),
    .io_in_b_valid(fb_io_in_b_valid),
    .io_in_ar_ready(fb_io_in_ar_ready),
    .io_in_ar_valid(fb_io_in_ar_valid),
    .io_in_ar_bits_addr(fb_io_in_ar_bits_addr),
    .io_in_r_ready(fb_io_in_r_ready),
    .io_in_r_valid(fb_io_in_r_valid),
    .io_in_r_bits_data(fb_io_in_r_bits_data)
  );
  FBHelper fbHelper ( // @[src/main/scala/device/AXI4VGA.scala 171:26]
    .clk(fbHelper_clk),
    .valid(fbHelper_valid),
    .pixel(fbHelper_pixel),
    .sync(fbHelper_sync)
  );
  GEN_w1_toggle #(.COVER_INDEX(10993)) toggle_10993 (
    .clock(toggle_10993_clock),
    .reset(toggle_10993_reset),
    .valid(toggle_10993_valid)
  );
  GEN_w11_toggle #(.COVER_INDEX(10994)) toggle_10994 (
    .clock(toggle_10994_clock),
    .reset(toggle_10994_reset),
    .valid(toggle_10994_valid)
  );
  GEN_w10_toggle #(.COVER_INDEX(11005)) toggle_11005 (
    .clock(toggle_11005_clock),
    .reset(toggle_11005_reset),
    .valid(toggle_11005_valid)
  );
  GEN_w17_toggle #(.COVER_INDEX(11015)) toggle_11015 (
    .clock(toggle_11015_clock),
    .reset(toggle_11015_reset),
    .valid(toggle_11015_valid)
  );
  GEN_w17_toggle #(.COVER_INDEX(11032)) toggle_11032 (
    .clock(toggle_11032_clock),
    .reset(toggle_11032_reset),
    .valid(toggle_11032_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(11049)) toggle_11049 (
    .clock(toggle_11049_clock),
    .reset(toggle_11049_reset),
    .valid(toggle_11049_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(11050)) toggle_11050 (
    .clock(toggle_11050_clock),
    .reset(toggle_11050_reset),
    .valid(toggle_11050_valid)
  );
  assign io_in_fb_aw_ready = fb_io_in_aw_ready; // @[src/main/scala/device/AXI4VGA.scala 130:15]
  assign io_in_fb_w_ready = fb_io_in_w_ready; // @[src/main/scala/device/AXI4VGA.scala 131:14]
  assign io_in_fb_b_valid = fb_io_in_b_valid; // @[src/main/scala/device/AXI4VGA.scala 132:14]
  assign io_in_fb_ar_ready = 1'h1; // @[src/main/scala/device/AXI4VGA.scala 133:21]
  assign io_in_fb_r_valid = io_in_fb_r_valid_r; // @[src/main/scala/device/AXI4VGA.scala 136:20]
  assign io_in_ctrl_aw_ready = ctrl_io_in_aw_ready; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign io_in_ctrl_w_ready = ctrl_io_in_w_ready; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign io_in_ctrl_b_valid = ctrl_io_in_b_valid; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign io_in_ctrl_ar_ready = ctrl_io_in_ar_ready; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign io_in_ctrl_r_valid = ctrl_io_in_r_valid; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign io_in_ctrl_r_bits_data = ctrl_io_in_r_bits_data; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign io_vga_valid = hInRange & vInRange; // @[src/main/scala/device/AXI4VGA.scala 148:28]
  assign ctrl_clock = clock;
  assign ctrl_reset = reset;
  assign ctrl_io_in_aw_valid = io_in_ctrl_aw_valid; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign ctrl_io_in_w_valid = io_in_ctrl_w_valid; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign ctrl_io_in_b_ready = io_in_ctrl_b_ready; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign ctrl_io_in_ar_valid = io_in_ctrl_ar_valid; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign ctrl_io_in_ar_bits_addr = io_in_ctrl_ar_bits_addr; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign ctrl_io_in_r_ready = io_in_ctrl_r_ready; // @[src/main/scala/device/AXI4VGA.scala 126:14]
  assign fb_clock = clock;
  assign fb_reset = reset;
  assign fb_io_in_aw_valid = io_in_fb_aw_valid; // @[src/main/scala/device/AXI4VGA.scala 130:15]
  assign fb_io_in_aw_bits_addr = io_in_fb_aw_bits_addr; // @[src/main/scala/device/AXI4VGA.scala 130:15]
  assign fb_io_in_w_valid = io_in_fb_w_valid; // @[src/main/scala/device/AXI4VGA.scala 131:14]
  assign fb_io_in_w_bits_data = io_in_fb_w_bits_data; // @[src/main/scala/device/AXI4VGA.scala 131:14]
  assign fb_io_in_w_bits_strb = io_in_fb_w_bits_strb; // @[src/main/scala/device/AXI4VGA.scala 131:14]
  assign fb_io_in_b_ready = io_in_fb_b_ready; // @[src/main/scala/device/AXI4VGA.scala 132:14]
  assign fb_io_in_ar_valid = fb_io_in_ar_valid_REG & hCounterIs2; // @[src/main/scala/device/AXI4VGA.scala 162:43]
  assign fb_io_in_ar_bits_addr = {{13'd0}, _fb_io_in_ar_bits_addr_T_1}; // @[src/main/scala/device/AXI4VGA.scala 161:25]
  assign fb_io_in_r_ready = 1'h1; // @[src/main/scala/device/AXI4VGA.scala 164:20]
  assign fbHelper_clk = clock; // @[src/main/scala/device/AXI4VGA.scala 172:21]
  assign fbHelper_valid = io_vga_valid; // @[src/main/scala/device/AXI4VGA.scala 173:23]
  assign fbHelper_pixel = hCounter[1] ? _GEN_14[63:32] : _GEN_14[31:0]; // @[src/main/scala/device/AXI4VGA.scala 167:23]
  assign fbHelper_sync = ctrl_io_extra_sync; // @[src/main/scala/device/AXI4VGA.scala 175:22]
  assign toggle_10993_clock = clock;
  assign toggle_10993_reset = reset;
  assign toggle_10993_valid = io_in_fb_r_valid_r ^ toggle_10993_valid_reg;
  assign toggle_10994_clock = clock;
  assign toggle_10994_reset = reset;
  assign toggle_10994_valid = hCounter ^ toggle_10994_valid_reg;
  assign toggle_11005_clock = clock;
  assign toggle_11005_reset = reset;
  assign toggle_11005_valid = vCounter ^ toggle_11005_valid_reg;
  assign toggle_11015_clock = clock;
  assign toggle_11015_reset = reset;
  assign toggle_11015_valid = fbPixelAddrV0 ^ toggle_11015_valid_reg;
  assign toggle_11032_clock = clock;
  assign toggle_11032_reset = reset;
  assign toggle_11032_valid = fbPixelAddrV1 ^ toggle_11032_valid_reg;
  assign toggle_11049_clock = clock;
  assign toggle_11049_reset = reset;
  assign toggle_11049_valid = fb_io_in_ar_valid_REG ^ toggle_11049_valid_reg;
  assign toggle_11050_clock = clock;
  assign toggle_11050_reset = reset;
  assign toggle_11050_valid = data_r ^ toggle_11050_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_fb_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_fb_r_valid_r <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      hCounter <= 11'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (wrap_wrap) begin // @[src/main/scala/chisel3/util/Counter.scala 87:20]
      hCounter <= 11'h0; // @[src/main/scala/chisel3/util/Counter.scala 87:28]
    end else begin
      hCounter <= _wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      vCounter <= 10'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (wrap_wrap) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      if (wrap_wrap_1) begin // @[src/main/scala/chisel3/util/Counter.scala 87:20]
        vCounter <= 10'h0; // @[src/main/scala/chisel3/util/Counter.scala 87:28]
      end else begin
        vCounter <= _wrap_value_T_3; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
      end
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      fbPixelAddrV0 <= 17'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_fbPixelAddrV0_T_1) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      if (fbPixelAddrV0_wrap_wrap) begin // @[src/main/scala/chisel3/util/Counter.scala 87:20]
        fbPixelAddrV0 <= 17'h0; // @[src/main/scala/chisel3/util/Counter.scala 87:28]
      end else begin
        fbPixelAddrV0 <= _fbPixelAddrV0_wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
      end
    end
    if (reset) begin // @[src/main/scala/chisel3/util/Counter.scala 61:40]
      fbPixelAddrV1 <= 17'h0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end else if (_fbPixelAddrV1_T) begin // @[src/main/scala/chisel3/util/Counter.scala 118:16]
      if (fbPixelAddrV1_wrap_wrap) begin // @[src/main/scala/chisel3/util/Counter.scala 87:20]
        fbPixelAddrV1 <= 17'h0; // @[src/main/scala/chisel3/util/Counter.scala 87:28]
      end else begin
        fbPixelAddrV1 <= _fbPixelAddrV1_wrap_value_T_1; // @[src/main/scala/chisel3/util/Counter.scala 77:15]
      end
    end
    fb_io_in_ar_valid_REG <= _nextPixel_T_2 & vInRange & hCounterIsOdd; // @[src/main/scala/device/AXI4VGA.scala 155:78]
    if (reset) begin // @[src/main/scala/utils/Hold.scala 23:65]
      data_r <= 64'h0; // @[src/main/scala/utils/Hold.scala 23:65]
    end else if (_data_T) begin // @[src/main/scala/utils/Hold.scala 23:65]
      data_r <= fb_io_in_r_bits_data; // @[src/main/scala/utils/Hold.scala 23:65]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    io_in_fb_r_valid_r_p <= io_in_fb_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_10993_valid_reg <= io_in_fb_r_valid_r;
    hCounter_p <= hCounter; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    toggle_10994_valid_reg <= hCounter;
    vCounter_p <= vCounter; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    toggle_11005_valid_reg <= vCounter;
    fbPixelAddrV0_p <= fbPixelAddrV0; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    toggle_11015_valid_reg <= fbPixelAddrV0;
    fbPixelAddrV1_p <= fbPixelAddrV1; // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    toggle_11032_valid_reg <= fbPixelAddrV1;
    fb_io_in_ar_valid_REG_p <= fb_io_in_ar_valid_REG; // @[src/main/scala/device/AXI4VGA.scala 162:31]
    toggle_11049_valid_reg <= fb_io_in_ar_valid_REG;
    data_r_p <= data_r; // @[src/main/scala/utils/Hold.scala 23:65]
    toggle_11050_valid_reg <= data_r;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_in_fb_r_valid_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  hCounter = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  vCounter = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  fbPixelAddrV0 = _RAND_3[16:0];
  _RAND_4 = {1{`RANDOM}};
  fbPixelAddrV1 = _RAND_4[16:0];
  _RAND_5 = {1{`RANDOM}};
  fb_io_in_ar_valid_REG = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  data_r = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  io_in_fb_r_valid_r_p = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  toggle_10993_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  hCounter_p = _RAND_9[10:0];
  _RAND_10 = {1{`RANDOM}};
  toggle_10994_valid_reg = _RAND_10[10:0];
  _RAND_11 = {1{`RANDOM}};
  vCounter_p = _RAND_11[9:0];
  _RAND_12 = {1{`RANDOM}};
  toggle_11005_valid_reg = _RAND_12[9:0];
  _RAND_13 = {1{`RANDOM}};
  fbPixelAddrV0_p = _RAND_13[16:0];
  _RAND_14 = {1{`RANDOM}};
  toggle_11015_valid_reg = _RAND_14[16:0];
  _RAND_15 = {1{`RANDOM}};
  fbPixelAddrV1_p = _RAND_15[16:0];
  _RAND_16 = {1{`RANDOM}};
  toggle_11032_valid_reg = _RAND_16[16:0];
  _RAND_17 = {1{`RANDOM}};
  fb_io_in_ar_valid_REG_p = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  toggle_11049_valid_reg = _RAND_18[0:0];
  _RAND_19 = {2{`RANDOM}};
  data_r_p = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  toggle_11050_valid_reg = _RAND_20[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(io_in_fb_r_valid_r_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(hCounter_t[0]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(hCounter_t[1]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(hCounter_t[2]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(hCounter_t[3]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(hCounter_t[4]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(hCounter_t[5]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(hCounter_t[6]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(hCounter_t[7]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(hCounter_t[8]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(hCounter_t[9]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(hCounter_t[10]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(vCounter_t[0]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(vCounter_t[1]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(vCounter_t[2]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(vCounter_t[3]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(vCounter_t[4]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(vCounter_t[5]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(vCounter_t[6]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(vCounter_t[7]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(vCounter_t[8]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(vCounter_t[9]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV0_t[0]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV0_t[1]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV0_t[2]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV0_t[3]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV0_t[4]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV0_t[5]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV0_t[6]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV0_t[7]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV0_t[8]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV0_t[9]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV0_t[10]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV0_t[11]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV0_t[12]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV0_t[13]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV0_t[14]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV0_t[15]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV0_t[16]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV1_t[0]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV1_t[1]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV1_t[2]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV1_t[3]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV1_t[4]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV1_t[5]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV1_t[6]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV1_t[7]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV1_t[8]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV1_t[9]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV1_t[10]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV1_t[11]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV1_t[12]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV1_t[13]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV1_t[14]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV1_t[15]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fbPixelAddrV1_t[16]); // @[src/main/scala/chisel3/util/Counter.scala 61:40]
    end
    //
    if (enToggle_past) begin
      cover(fb_io_in_ar_valid_REG_t); // @[src/main/scala/device/AXI4VGA.scala 162:31]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[0]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[1]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[2]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[3]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[4]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[5]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[6]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[7]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[8]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[9]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[10]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[11]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[12]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[13]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[14]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[15]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[16]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[17]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[18]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[19]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[20]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[21]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[22]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[23]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[24]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[25]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[26]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[27]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[28]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[29]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[30]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[31]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[32]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[33]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[34]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[35]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[36]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[37]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[38]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[39]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[40]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[41]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[42]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[43]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[44]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[45]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[46]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[47]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[48]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[49]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[50]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[51]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[52]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[53]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[54]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[55]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[56]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[57]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[58]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[59]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[60]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[61]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[62]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
    //
    if (enToggle_past) begin
      cover(data_r_t[63]); // @[src/main/scala/utils/Hold.scala 23:65]
    end
  end
endmodule
module AXI4Flash(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire  _r_busy_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _r_busy_T_1 = io_in_r_ready & io_in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _r_busy_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_2 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io_in_b_ready & io_in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _w_busy_T | _GEN_4; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _rdata_T = 11'h0 == io_in_ar_bits_addr[12:2]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_1 = 11'h1 == io_in_ar_bits_addr[12:2]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_2 = 11'h2 == io_in_ar_bits_addr[12:2]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [20:0] _rdata_T_3 = _rdata_T ? 21'h10029b : 21'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [24:0] _rdata_T_4 = _rdata_T_1 ? 25'h1f29293 : 25'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [17:0] _rdata_T_5 = _rdata_T_2 ? 18'h28067 : 18'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [24:0] _GEN_15 = {{4'd0}, _rdata_T_3}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [24:0] _rdata_T_6 = _GEN_15 | _rdata_T_4; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [24:0] _GEN_16 = {{7'd0}, _rdata_T_5}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [24:0] _rdata_T_7 = _rdata_T_6 | _GEN_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [63:0] rdata = {{39'd0}, _rdata_T_7}; // @[src/main/scala/device/AXI4Flash.scala 37:19 src/main/scala/utils/RegMap.scala 30:11]
  reg [63:0] io_in_r_bits_data_REG; // @[src/main/scala/device/AXI4Flash.scala 41:38]
  reg [63:0] io_in_r_bits_data_r; // @[src/main/scala/device/AXI4Flash.scala 41:30]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  r_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  r_busy_t = r_busy ^ r_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_11114_clock;
  wire  toggle_11114_reset;
  wire  toggle_11114_valid;
  reg  toggle_11114_valid_reg;
  reg  ren_REG_p; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  ren_REG_t = ren_REG ^ ren_REG_p; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  toggle_11115_clock;
  wire  toggle_11115_reset;
  wire  toggle_11115_valid;
  reg  toggle_11115_valid_reg;
  reg  io_in_r_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  io_in_r_valid_r_t = io_in_r_valid_r ^ io_in_r_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_11116_clock;
  wire  toggle_11116_reset;
  wire  toggle_11116_valid;
  reg  toggle_11116_valid_reg;
  reg  w_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  w_busy_t = w_busy ^ w_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_11117_clock;
  wire  toggle_11117_reset;
  wire  toggle_11117_valid;
  reg  toggle_11117_valid_reg;
  reg  io_in_b_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  io_in_b_valid_r_t = io_in_b_valid_r ^ io_in_b_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_11118_clock;
  wire  toggle_11118_reset;
  wire  toggle_11118_valid;
  reg  toggle_11118_valid_reg;
  reg [63:0] io_in_r_bits_data_REG_p; // @[src/main/scala/device/AXI4Flash.scala 41:38]
  wire [63:0] io_in_r_bits_data_REG_t = io_in_r_bits_data_REG ^ io_in_r_bits_data_REG_p; // @[src/main/scala/device/AXI4Flash.scala 41:38]
  wire  toggle_11119_clock;
  wire  toggle_11119_reset;
  wire [63:0] toggle_11119_valid;
  reg [63:0] toggle_11119_valid_reg;
  reg [63:0] io_in_r_bits_data_r_p; // @[src/main/scala/device/AXI4Flash.scala 41:30]
  wire [63:0] io_in_r_bits_data_r_t = io_in_r_bits_data_r ^ io_in_r_bits_data_r_p; // @[src/main/scala/device/AXI4Flash.scala 41:30]
  wire  toggle_11183_clock;
  wire  toggle_11183_reset;
  wire [63:0] toggle_11183_valid;
  reg [63:0] toggle_11183_valid_reg;
  GEN_w1_toggle #(.COVER_INDEX(11114)) toggle_11114 (
    .clock(toggle_11114_clock),
    .reset(toggle_11114_reset),
    .valid(toggle_11114_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(11115)) toggle_11115 (
    .clock(toggle_11115_clock),
    .reset(toggle_11115_reset),
    .valid(toggle_11115_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(11116)) toggle_11116 (
    .clock(toggle_11116_clock),
    .reset(toggle_11116_reset),
    .valid(toggle_11116_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(11117)) toggle_11117 (
    .clock(toggle_11117_clock),
    .reset(toggle_11117_reset),
    .valid(toggle_11117_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(11118)) toggle_11118 (
    .clock(toggle_11118_clock),
    .reset(toggle_11118_reset),
    .valid(toggle_11118_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(11119)) toggle_11119 (
    .clock(toggle_11119_clock),
    .reset(toggle_11119_reset),
    .valid(toggle_11119_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(11183)) toggle_11183 (
    .clock(toggle_11183_clock),
    .reset(toggle_11183_reset),
    .valid(toggle_11183_valid)
  );
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = io_in_r_bits_data_r; // @[src/main/scala/device/AXI4Flash.scala 41:18]
  assign toggle_11114_clock = clock;
  assign toggle_11114_reset = reset;
  assign toggle_11114_valid = r_busy ^ toggle_11114_valid_reg;
  assign toggle_11115_clock = clock;
  assign toggle_11115_reset = reset;
  assign toggle_11115_valid = ren_REG ^ toggle_11115_valid_reg;
  assign toggle_11116_clock = clock;
  assign toggle_11116_reset = reset;
  assign toggle_11116_valid = io_in_r_valid_r ^ toggle_11116_valid_reg;
  assign toggle_11117_clock = clock;
  assign toggle_11117_reset = reset;
  assign toggle_11117_valid = w_busy ^ toggle_11117_valid_reg;
  assign toggle_11118_clock = clock;
  assign toggle_11118_reset = reset;
  assign toggle_11118_valid = io_in_b_valid_r ^ toggle_11118_valid_reg;
  assign toggle_11119_clock = clock;
  assign toggle_11119_reset = reset;
  assign toggle_11119_valid = io_in_r_bits_data_REG ^ toggle_11119_valid_reg;
  assign toggle_11183_clock = clock;
  assign toggle_11183_reset = reset;
  assign toggle_11183_valid = io_in_r_bits_data_r ^ toggle_11183_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
    io_in_r_bits_data_REG <= {rdata[31:0],rdata[31:0]}; // @[src/main/scala/device/AXI4Flash.scala 41:43]
    if (ren_REG) begin // @[src/main/scala/device/AXI4Flash.scala 41:30]
      io_in_r_bits_data_r <= io_in_r_bits_data_REG; // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    r_busy_p <= r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_11114_valid_reg <= r_busy;
    ren_REG_p <= ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    toggle_11115_valid_reg <= ren_REG;
    io_in_r_valid_r_p <= io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_11116_valid_reg <= io_in_r_valid_r;
    w_busy_p <= w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_11117_valid_reg <= w_busy;
    io_in_b_valid_r_p <= io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_11118_valid_reg <= io_in_b_valid_r;
    io_in_r_bits_data_REG_p <= io_in_r_bits_data_REG; // @[src/main/scala/device/AXI4Flash.scala 41:38]
    toggle_11119_valid_reg <= io_in_r_bits_data_REG;
    io_in_r_bits_data_r_p <= io_in_r_bits_data_r; // @[src/main/scala/device/AXI4Flash.scala 41:30]
    toggle_11183_valid_reg <= io_in_r_bits_data_r;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  io_in_r_bits_data_REG = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  io_in_r_bits_data_r = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  r_busy_p = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  toggle_11114_valid_reg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  ren_REG_p = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  toggle_11115_valid_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  io_in_r_valid_r_p = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  toggle_11116_valid_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  w_busy_p = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  toggle_11117_valid_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  io_in_b_valid_r_p = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  toggle_11118_valid_reg = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  io_in_r_bits_data_REG_p = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  toggle_11119_valid_reg = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  io_in_r_bits_data_r_p = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  toggle_11183_valid_reg = _RAND_20[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(r_busy_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(ren_REG_t); // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_valid_r_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(w_busy_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(io_in_b_valid_r_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[0]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[1]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[2]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[3]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[4]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[5]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[6]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[7]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[8]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[9]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[10]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[11]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[12]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[13]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[14]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[15]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[16]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[17]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[18]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[19]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[20]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[21]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[22]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[23]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[24]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[25]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[26]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[27]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[28]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[29]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[30]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[31]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[32]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[33]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[34]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[35]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[36]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[37]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[38]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[39]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[40]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[41]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[42]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[43]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[44]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[45]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[46]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[47]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[48]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[49]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[50]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[51]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[52]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[53]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[54]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[55]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[56]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[57]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[58]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[59]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[60]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[61]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[62]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[63]); // @[src/main/scala/device/AXI4Flash.scala 41:38]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[0]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[1]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[2]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[3]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[4]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[5]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[6]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[7]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[8]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[9]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[10]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[11]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[12]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[13]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[14]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[15]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[16]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[17]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[18]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[19]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[20]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[21]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[22]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[23]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[24]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[25]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[26]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[27]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[28]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[29]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[30]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[31]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[32]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[33]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[34]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[35]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[36]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[37]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[38]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[39]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[40]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[41]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[42]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[43]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[44]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[45]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[46]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[47]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[48]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[49]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[50]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[51]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[52]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[53]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[54]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[55]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[56]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[57]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[58]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[59]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[60]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[61]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[62]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[63]); // @[src/main/scala/device/AXI4Flash.scala 41:30]
    end
  end
endmodule
module AXI4DummySD(
  input         clock,
  input         reset,
  output        io_in_aw_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_aw_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_aw_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_w_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_w_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [63:0] io_in_w_bits_data, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [7:0]  io_in_w_bits_strb, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_b_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_b_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_ar_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_ar_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input  [31:0] io_in_ar_bits_addr, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  input         io_in_r_ready, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output        io_in_r_valid, // @[src/main/scala/device/AXI4Slave.scala 28:14]
  output [63:0] io_in_r_bits_data // @[src/main/scala/device/AXI4Slave.scala 28:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
`endif // RANDOMIZE_REG_INIT
  wire  sdHelper_clk; // @[src/main/scala/device/AXI4DummySD.scala 114:24]
  wire  sdHelper_ren; // @[src/main/scala/device/AXI4DummySD.scala 114:24]
  wire [31:0] sdHelper_data; // @[src/main/scala/device/AXI4DummySD.scala 114:24]
  wire  sdHelper_setAddr; // @[src/main/scala/device/AXI4DummySD.scala 114:24]
  wire [31:0] sdHelper_addr; // @[src/main/scala/device/AXI4DummySD.scala 114:24]
  wire  _r_busy_T = io_in_ar_ready & io_in_ar_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _r_busy_T_1 = io_in_r_ready & io_in_r_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _r_busy_T_1 ? 1'h0 : r_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_1 = _r_busy_T | _GEN_0; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg  ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  _io_in_r_valid_T_2 = ren_REG & (_r_busy_T | r_busy); // @[src/main/scala/device/AXI4Slave.scala 74:35]
  reg  io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_2 = _r_busy_T_1 ? 1'h0 : io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_3 = _io_in_r_valid_T_2 | _GEN_2; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _w_busy_T = io_in_aw_ready & io_in_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  wire  _w_busy_T_1 = io_in_b_ready & io_in_b_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_4 = _w_busy_T_1 ? 1'h0 : w_busy; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_5 = _w_busy_T | _GEN_4; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  wire  _io_in_b_valid_T = io_in_w_ready & io_in_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_6 = _w_busy_T_1 ? 1'h0 : io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 26:19 24:20 26:23]
  wire  _GEN_7 = _io_in_b_valid_T | _GEN_6; // @[src/main/scala/utils/StopWatch.scala 27:{20,24}]
  reg [31:0] regs_0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_1; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_4; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_5; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_6; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_7; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_8; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_15; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  reg [31:0] regs_20; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire [3:0] strb = io_in_aw_bits_addr[2] ? io_in_w_bits_strb[7:4] : io_in_w_bits_strb[3:0]; // @[src/main/scala/device/AXI4DummySD.scala 138:22]
  wire [7:0] _T_8 = strb[0] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_9 = strb[1] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_10 = strb[2] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [7:0] _T_11 = strb[3] ? 8'hff : 8'h0; // @[src/main/scala/utils/BitUtils.scala 27:46]
  wire [31:0] _T_12 = {_T_11,_T_10,_T_9,_T_8}; // @[src/main/scala/utils/BitUtils.scala 27:27]
  wire  _rdata_T = 13'h0 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_1 = 13'h38 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_2 = 13'h18 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_3 = 13'h34 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_4 = 13'h14 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_5 = 13'h1c == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_6 = 13'h50 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_7 = 13'h10 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_8 = 13'h4 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_9 = 13'h20 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire  _rdata_T_10 = 13'h40 == io_in_ar_bits_addr[12:0]; // @[src/main/scala/utils/LookupTree.scala 24:34]
  wire [31:0] _rdata_T_11 = _rdata_T ? regs_0 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_12 = _rdata_T_1 ? regs_15 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_13 = _rdata_T_2 ? regs_6 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [7:0] _rdata_T_14 = _rdata_T_3 ? 8'h80 : 8'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_15 = _rdata_T_4 ? regs_5 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_16 = _rdata_T_5 ? regs_7 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_17 = _rdata_T_6 ? regs_20 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_18 = _rdata_T_7 ? regs_4 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_19 = _rdata_T_8 ? regs_1 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_20 = _rdata_T_9 ? regs_8 : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_21 = _rdata_T_10 ? sdHelper_data : 32'h0; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_22 = _rdata_T_11 | _rdata_T_12; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_23 = _rdata_T_22 | _rdata_T_13; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _GEN_53 = {{24'd0}, _rdata_T_14}; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_24 = _rdata_T_23 | _GEN_53; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_25 = _rdata_T_24 | _rdata_T_15; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_26 = _rdata_T_25 | _rdata_T_16; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_27 = _rdata_T_26 | _rdata_T_17; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_28 = _rdata_T_27 | _rdata_T_18; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_29 = _rdata_T_28 | _rdata_T_19; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_30 = _rdata_T_29 | _rdata_T_20; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _rdata_T_31 = _rdata_T_30 | _rdata_T_21; // @[src/main/scala/chisel3/util/Mux.scala 30:73]
  wire [31:0] _regs_0_T = io_in_w_bits_data[31:0] & _T_12; // @[src/main/scala/utils/BitUtils.scala 34:14]
  wire [31:0] _regs_0_T_1 = ~_T_12; // @[src/main/scala/utils/BitUtils.scala 34:39]
  wire [31:0] _regs_0_T_2 = regs_0 & _regs_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _regs_0_T_3 = _regs_0_T | _regs_0_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [5:0] regs_0_cmd = _regs_0_T_3[5:0]; // @[src/main/scala/device/AXI4DummySD.scala 84:20]
  wire [31:0] _GEN_9 = 6'hd == regs_0_cmd ? 32'h0 : regs_4; // @[src/main/scala/device/AXI4DummySD.scala 85:18 102:22 72:43]
  wire [31:0] _GEN_10 = 6'hd == regs_0_cmd ? 32'h0 : regs_5; // @[src/main/scala/device/AXI4DummySD.scala 85:18 103:22 72:43]
  wire [31:0] _GEN_11 = 6'hd == regs_0_cmd ? 32'h0 : regs_6; // @[src/main/scala/device/AXI4DummySD.scala 85:18 104:22 72:43]
  wire [31:0] _GEN_12 = 6'hd == regs_0_cmd ? 32'h0 : regs_7; // @[src/main/scala/device/AXI4DummySD.scala 85:18 105:22 72:43]
  wire  _GEN_13 = 6'hd == regs_0_cmd ? 1'h0 : 6'h12 == regs_0_cmd; // @[src/main/scala/device/AXI4DummySD.scala 85:18 81:25]
  wire [31:0] _GEN_14 = 6'h9 == regs_0_cmd ? 32'h92404001 : _GEN_9; // @[src/main/scala/device/AXI4DummySD.scala 85:18 96:22]
  wire [31:0] _GEN_15 = 6'h9 == regs_0_cmd ? 32'hd24b97e3 : _GEN_10; // @[src/main/scala/device/AXI4DummySD.scala 85:18 97:22]
  wire [31:0] _GEN_16 = 6'h9 == regs_0_cmd ? 32'hf5f803f : _GEN_11; // @[src/main/scala/device/AXI4DummySD.scala 85:18 98:22]
  wire [31:0] _GEN_17 = 6'h9 == regs_0_cmd ? 32'h8c26012a : _GEN_12; // @[src/main/scala/device/AXI4DummySD.scala 85:18 99:22]
  wire  _GEN_18 = 6'h9 == regs_0_cmd ? 1'h0 : _GEN_13; // @[src/main/scala/device/AXI4DummySD.scala 85:18 81:25]
  wire  _GEN_23 = 6'h2 == regs_0_cmd ? 1'h0 : _GEN_18; // @[src/main/scala/device/AXI4DummySD.scala 85:18 81:25]
  wire  _GEN_28 = 6'h1 == regs_0_cmd ? 1'h0 : _GEN_23; // @[src/main/scala/device/AXI4DummySD.scala 85:18 81:25]
  wire [31:0] _regs_15_T_2 = regs_15 & _regs_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _regs_15_T_3 = _regs_0_T | _regs_15_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _regs_20_T_2 = regs_20 & _regs_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _regs_20_T_3 = _regs_0_T | _regs_20_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _regs_1_T_2 = regs_1 & _regs_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _regs_1_T_3 = _regs_0_T | _regs_1_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [31:0] _regs_8_T_2 = regs_8 & _regs_0_T_1; // @[src/main/scala/utils/BitUtils.scala 34:37]
  wire [31:0] _regs_8_T_3 = _regs_0_T | _regs_8_T_2; // @[src/main/scala/utils/BitUtils.scala 34:26]
  wire [63:0] rdata = {{32'd0}, _rdata_T_31}; // @[src/main/scala/device/AXI4DummySD.scala 139:19 src/main/scala/utils/RegMap.scala 30:11]
  reg [63:0] io_in_r_bits_data_REG; // @[src/main/scala/device/AXI4DummySD.scala 144:44]
  reg [63:0] io_in_r_bits_data_r; // @[src/main/scala/device/AXI4DummySD.scala 144:36]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  r_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  r_busy_t = r_busy ^ r_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_11247_clock;
  wire  toggle_11247_reset;
  wire  toggle_11247_valid;
  reg  toggle_11247_valid_reg;
  reg  ren_REG_p; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  ren_REG_t = ren_REG ^ ren_REG_p; // @[src/main/scala/device/AXI4Slave.scala 73:17]
  wire  toggle_11248_clock;
  wire  toggle_11248_reset;
  wire  toggle_11248_valid;
  reg  toggle_11248_valid_reg;
  reg  io_in_r_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  io_in_r_valid_r_t = io_in_r_valid_r ^ io_in_r_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_11249_clock;
  wire  toggle_11249_reset;
  wire  toggle_11249_valid;
  reg  toggle_11249_valid_reg;
  reg  w_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  w_busy_t = w_busy ^ w_busy_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_11250_clock;
  wire  toggle_11250_reset;
  wire  toggle_11250_valid;
  reg  toggle_11250_valid_reg;
  reg  io_in_b_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  io_in_b_valid_r_t = io_in_b_valid_r ^ io_in_b_valid_r_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_11251_clock;
  wire  toggle_11251_reset;
  wire  toggle_11251_valid;
  reg  toggle_11251_valid_reg;
  reg [31:0] regs_0_p; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire [31:0] regs_0_t = regs_0 ^ regs_0_p; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire  toggle_11252_clock;
  wire  toggle_11252_reset;
  wire [31:0] toggle_11252_valid;
  reg [31:0] toggle_11252_valid_reg;
  reg [31:0] regs_1_p; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire [31:0] regs_1_t = regs_1 ^ regs_1_p; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire  toggle_11284_clock;
  wire  toggle_11284_reset;
  wire [31:0] toggle_11284_valid;
  reg [31:0] toggle_11284_valid_reg;
  reg [31:0] regs_4_p; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire [31:0] regs_4_t = regs_4 ^ regs_4_p; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire  toggle_11316_clock;
  wire  toggle_11316_reset;
  wire [31:0] toggle_11316_valid;
  reg [31:0] toggle_11316_valid_reg;
  reg [31:0] regs_5_p; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire [31:0] regs_5_t = regs_5 ^ regs_5_p; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire  toggle_11348_clock;
  wire  toggle_11348_reset;
  wire [31:0] toggle_11348_valid;
  reg [31:0] toggle_11348_valid_reg;
  reg [31:0] regs_6_p; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire [31:0] regs_6_t = regs_6 ^ regs_6_p; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire  toggle_11380_clock;
  wire  toggle_11380_reset;
  wire [31:0] toggle_11380_valid;
  reg [31:0] toggle_11380_valid_reg;
  reg [31:0] regs_7_p; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire [31:0] regs_7_t = regs_7 ^ regs_7_p; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire  toggle_11412_clock;
  wire  toggle_11412_reset;
  wire [31:0] toggle_11412_valid;
  reg [31:0] toggle_11412_valid_reg;
  reg [31:0] regs_8_p; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire [31:0] regs_8_t = regs_8 ^ regs_8_p; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire  toggle_11444_clock;
  wire  toggle_11444_reset;
  wire [31:0] toggle_11444_valid;
  reg [31:0] toggle_11444_valid_reg;
  reg [31:0] regs_15_p; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire [31:0] regs_15_t = regs_15 ^ regs_15_p; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire  toggle_11476_clock;
  wire  toggle_11476_reset;
  wire [31:0] toggle_11476_valid;
  reg [31:0] toggle_11476_valid_reg;
  reg [31:0] regs_20_p; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire [31:0] regs_20_t = regs_20 ^ regs_20_p; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
  wire  toggle_11508_clock;
  wire  toggle_11508_reset;
  wire [31:0] toggle_11508_valid;
  reg [31:0] toggle_11508_valid_reg;
  reg [63:0] io_in_r_bits_data_REG_p; // @[src/main/scala/device/AXI4DummySD.scala 144:44]
  wire [63:0] io_in_r_bits_data_REG_t = io_in_r_bits_data_REG ^ io_in_r_bits_data_REG_p; // @[src/main/scala/device/AXI4DummySD.scala 144:44]
  wire  toggle_11540_clock;
  wire  toggle_11540_reset;
  wire [63:0] toggle_11540_valid;
  reg [63:0] toggle_11540_valid_reg;
  reg [63:0] io_in_r_bits_data_r_p; // @[src/main/scala/device/AXI4DummySD.scala 144:36]
  wire [63:0] io_in_r_bits_data_r_t = io_in_r_bits_data_r ^ io_in_r_bits_data_r_p; // @[src/main/scala/device/AXI4DummySD.scala 144:36]
  wire  toggle_11604_clock;
  wire  toggle_11604_reset;
  wire [63:0] toggle_11604_valid;
  reg [63:0] toggle_11604_valid_reg;
  SDHelper sdHelper ( // @[src/main/scala/device/AXI4DummySD.scala 114:24]
    .clk(sdHelper_clk),
    .ren(sdHelper_ren),
    .data(sdHelper_data),
    .setAddr(sdHelper_setAddr),
    .addr(sdHelper_addr)
  );
  GEN_w1_toggle #(.COVER_INDEX(11247)) toggle_11247 (
    .clock(toggle_11247_clock),
    .reset(toggle_11247_reset),
    .valid(toggle_11247_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(11248)) toggle_11248 (
    .clock(toggle_11248_clock),
    .reset(toggle_11248_reset),
    .valid(toggle_11248_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(11249)) toggle_11249 (
    .clock(toggle_11249_clock),
    .reset(toggle_11249_reset),
    .valid(toggle_11249_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(11250)) toggle_11250 (
    .clock(toggle_11250_clock),
    .reset(toggle_11250_reset),
    .valid(toggle_11250_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(11251)) toggle_11251 (
    .clock(toggle_11251_clock),
    .reset(toggle_11251_reset),
    .valid(toggle_11251_valid)
  );
  GEN_w32_toggle #(.COVER_INDEX(11252)) toggle_11252 (
    .clock(toggle_11252_clock),
    .reset(toggle_11252_reset),
    .valid(toggle_11252_valid)
  );
  GEN_w32_toggle #(.COVER_INDEX(11284)) toggle_11284 (
    .clock(toggle_11284_clock),
    .reset(toggle_11284_reset),
    .valid(toggle_11284_valid)
  );
  GEN_w32_toggle #(.COVER_INDEX(11316)) toggle_11316 (
    .clock(toggle_11316_clock),
    .reset(toggle_11316_reset),
    .valid(toggle_11316_valid)
  );
  GEN_w32_toggle #(.COVER_INDEX(11348)) toggle_11348 (
    .clock(toggle_11348_clock),
    .reset(toggle_11348_reset),
    .valid(toggle_11348_valid)
  );
  GEN_w32_toggle #(.COVER_INDEX(11380)) toggle_11380 (
    .clock(toggle_11380_clock),
    .reset(toggle_11380_reset),
    .valid(toggle_11380_valid)
  );
  GEN_w32_toggle #(.COVER_INDEX(11412)) toggle_11412 (
    .clock(toggle_11412_clock),
    .reset(toggle_11412_reset),
    .valid(toggle_11412_valid)
  );
  GEN_w32_toggle #(.COVER_INDEX(11444)) toggle_11444 (
    .clock(toggle_11444_clock),
    .reset(toggle_11444_reset),
    .valid(toggle_11444_valid)
  );
  GEN_w32_toggle #(.COVER_INDEX(11476)) toggle_11476 (
    .clock(toggle_11476_clock),
    .reset(toggle_11476_reset),
    .valid(toggle_11476_valid)
  );
  GEN_w32_toggle #(.COVER_INDEX(11508)) toggle_11508 (
    .clock(toggle_11508_clock),
    .reset(toggle_11508_reset),
    .valid(toggle_11508_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(11540)) toggle_11540 (
    .clock(toggle_11540_clock),
    .reset(toggle_11540_reset),
    .valid(toggle_11540_valid)
  );
  GEN_w64_toggle #(.COVER_INDEX(11604)) toggle_11604 (
    .clock(toggle_11604_clock),
    .reset(toggle_11604_reset),
    .valid(toggle_11604_valid)
  );
  assign io_in_aw_ready = ~w_busy; // @[src/main/scala/device/AXI4Slave.scala 94:18]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[src/main/scala/device/AXI4Slave.scala 95:30]
  assign io_in_b_valid = io_in_b_valid_r; // @[src/main/scala/device/AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | ~r_busy; // @[src/main/scala/device/AXI4Slave.scala 71:29]
  assign io_in_r_valid = io_in_r_valid_r; // @[src/main/scala/device/AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = io_in_r_bits_data_r; // @[src/main/scala/device/AXI4DummySD.scala 143:18]
  assign sdHelper_clk = clock; // @[src/main/scala/device/AXI4DummySD.scala 115:19]
  assign sdHelper_ren = io_in_ar_bits_addr[12:0] == 13'h40 & _r_busy_T; // @[src/main/scala/device/AXI4DummySD.scala 116:51]
  assign sdHelper_setAddr = _io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h0 & _GEN_28; // @[src/main/scala/utils/RegMap.scala 32:48 src/main/scala/device/AXI4DummySD.scala 81:25]
  assign sdHelper_addr = regs_1; // @[src/main/scala/device/AXI4DummySD.scala 118:20]
  assign toggle_11247_clock = clock;
  assign toggle_11247_reset = reset;
  assign toggle_11247_valid = r_busy ^ toggle_11247_valid_reg;
  assign toggle_11248_clock = clock;
  assign toggle_11248_reset = reset;
  assign toggle_11248_valid = ren_REG ^ toggle_11248_valid_reg;
  assign toggle_11249_clock = clock;
  assign toggle_11249_reset = reset;
  assign toggle_11249_valid = io_in_r_valid_r ^ toggle_11249_valid_reg;
  assign toggle_11250_clock = clock;
  assign toggle_11250_reset = reset;
  assign toggle_11250_valid = w_busy ^ toggle_11250_valid_reg;
  assign toggle_11251_clock = clock;
  assign toggle_11251_reset = reset;
  assign toggle_11251_valid = io_in_b_valid_r ^ toggle_11251_valid_reg;
  assign toggle_11252_clock = clock;
  assign toggle_11252_reset = reset;
  assign toggle_11252_valid = regs_0 ^ toggle_11252_valid_reg;
  assign toggle_11284_clock = clock;
  assign toggle_11284_reset = reset;
  assign toggle_11284_valid = regs_1 ^ toggle_11284_valid_reg;
  assign toggle_11316_clock = clock;
  assign toggle_11316_reset = reset;
  assign toggle_11316_valid = regs_4 ^ toggle_11316_valid_reg;
  assign toggle_11348_clock = clock;
  assign toggle_11348_reset = reset;
  assign toggle_11348_valid = regs_5 ^ toggle_11348_valid_reg;
  assign toggle_11380_clock = clock;
  assign toggle_11380_reset = reset;
  assign toggle_11380_valid = regs_6 ^ toggle_11380_valid_reg;
  assign toggle_11412_clock = clock;
  assign toggle_11412_reset = reset;
  assign toggle_11412_valid = regs_7 ^ toggle_11412_valid_reg;
  assign toggle_11444_clock = clock;
  assign toggle_11444_reset = reset;
  assign toggle_11444_valid = regs_8 ^ toggle_11444_valid_reg;
  assign toggle_11476_clock = clock;
  assign toggle_11476_reset = reset;
  assign toggle_11476_valid = regs_15 ^ toggle_11476_valid_reg;
  assign toggle_11508_clock = clock;
  assign toggle_11508_reset = reset;
  assign toggle_11508_valid = regs_20 ^ toggle_11508_valid_reg;
  assign toggle_11540_clock = clock;
  assign toggle_11540_reset = reset;
  assign toggle_11540_valid = io_in_r_bits_data_REG ^ toggle_11540_valid_reg;
  assign toggle_11604_clock = clock;
  assign toggle_11604_reset = reset;
  assign toggle_11604_valid = io_in_r_bits_data_r ^ toggle_11604_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[src/main/scala/device/AXI4Slave.scala 73:17]
      ren_REG <= 1'h0; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end else begin
      ren_REG <= _r_busy_T; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_r_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_r_valid_r <= _GEN_3;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      io_in_b_valid_r <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else begin
      io_in_b_valid_r <= _GEN_7;
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_0 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      regs_0 <= _regs_0_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_1 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h4) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      regs_1 <= _regs_1_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_4 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      if (6'h1 == regs_0_cmd) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
        regs_4 <= 32'h80ff8000; // @[src/main/scala/device/AXI4DummySD.scala 87:22]
      end else if (6'h2 == regs_0_cmd) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
        regs_4 <= 32'h1; // @[src/main/scala/device/AXI4DummySD.scala 90:22]
      end else begin
        regs_4 <= _GEN_14;
      end
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_5 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      if (!(6'h1 == regs_0_cmd)) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
        if (6'h2 == regs_0_cmd) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
          regs_5 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 91:22]
        end else begin
          regs_5 <= _GEN_15;
        end
      end
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_6 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      if (!(6'h1 == regs_0_cmd)) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
        if (6'h2 == regs_0_cmd) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
          regs_6 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 92:22]
        end else begin
          regs_6 <= _GEN_16;
        end
      end
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_7 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h0) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      if (!(6'h1 == regs_0_cmd)) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
        if (6'h2 == regs_0_cmd) begin // @[src/main/scala/device/AXI4DummySD.scala 85:18]
          regs_7 <= 32'h15000000; // @[src/main/scala/device/AXI4DummySD.scala 93:22]
        end else begin
          regs_7 <= _GEN_17;
        end
      end
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_8 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h20) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      regs_8 <= _regs_8_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_15 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h38) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      regs_15 <= _regs_15_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    if (reset) begin // @[src/main/scala/device/AXI4DummySD.scala 72:43]
      regs_20 <= 32'h0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end else if (_io_in_b_valid_T & io_in_aw_bits_addr[12:0] == 13'h50) begin // @[src/main/scala/utils/RegMap.scala 32:48]
      regs_20 <= _regs_20_T_3; // @[src/main/scala/utils/RegMap.scala 32:52]
    end
    io_in_r_bits_data_REG <= {rdata[31:0],rdata[31:0]}; // @[src/main/scala/device/AXI4DummySD.scala 144:49]
    if (ren_REG) begin // @[src/main/scala/device/AXI4DummySD.scala 144:36]
      io_in_r_bits_data_r <= io_in_r_bits_data_REG; // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    r_busy_p <= r_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_11247_valid_reg <= r_busy;
    ren_REG_p <= ren_REG; // @[src/main/scala/device/AXI4Slave.scala 73:17]
    toggle_11248_valid_reg <= ren_REG;
    io_in_r_valid_r_p <= io_in_r_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_11249_valid_reg <= io_in_r_valid_r;
    w_busy_p <= w_busy; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_11250_valid_reg <= w_busy;
    io_in_b_valid_r_p <= io_in_b_valid_r; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_11251_valid_reg <= io_in_b_valid_r;
    regs_0_p <= regs_0; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    toggle_11252_valid_reg <= regs_0;
    regs_1_p <= regs_1; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    toggle_11284_valid_reg <= regs_1;
    regs_4_p <= regs_4; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    toggle_11316_valid_reg <= regs_4;
    regs_5_p <= regs_5; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    toggle_11348_valid_reg <= regs_5;
    regs_6_p <= regs_6; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    toggle_11380_valid_reg <= regs_6;
    regs_7_p <= regs_7; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    toggle_11412_valid_reg <= regs_7;
    regs_8_p <= regs_8; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    toggle_11444_valid_reg <= regs_8;
    regs_15_p <= regs_15; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    toggle_11476_valid_reg <= regs_15;
    regs_20_p <= regs_20; // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    toggle_11508_valid_reg <= regs_20;
    io_in_r_bits_data_REG_p <= io_in_r_bits_data_REG; // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    toggle_11540_valid_reg <= io_in_r_bits_data_REG;
    io_in_r_bits_data_r_p <= io_in_r_bits_data_r; // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    toggle_11604_valid_reg <= io_in_r_bits_data_r;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_in_r_valid_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_in_b_valid_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  regs_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regs_1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regs_4 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regs_5 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regs_6 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regs_7 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regs_8 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regs_15 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  regs_20 = _RAND_13[31:0];
  _RAND_14 = {2{`RANDOM}};
  io_in_r_bits_data_REG = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  io_in_r_bits_data_r = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  r_busy_p = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  toggle_11247_valid_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  ren_REG_p = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  toggle_11248_valid_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  io_in_r_valid_r_p = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  toggle_11249_valid_reg = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  w_busy_p = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  toggle_11250_valid_reg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  io_in_b_valid_r_p = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  toggle_11251_valid_reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  regs_0_p = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  toggle_11252_valid_reg = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  regs_1_p = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  toggle_11284_valid_reg = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  regs_4_p = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  toggle_11316_valid_reg = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  regs_5_p = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  toggle_11348_valid_reg = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  regs_6_p = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  toggle_11380_valid_reg = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  regs_7_p = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  toggle_11412_valid_reg = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  regs_8_p = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  toggle_11444_valid_reg = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  regs_15_p = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  toggle_11476_valid_reg = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  regs_20_p = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  toggle_11508_valid_reg = _RAND_43[31:0];
  _RAND_44 = {2{`RANDOM}};
  io_in_r_bits_data_REG_p = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  toggle_11540_valid_reg = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  io_in_r_bits_data_r_p = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  toggle_11604_valid_reg = _RAND_47[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (enToggle_past) begin
      cover(r_busy_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(ren_REG_t); // @[src/main/scala/device/AXI4Slave.scala 73:17]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_valid_r_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(w_busy_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(io_in_b_valid_r_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[0]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[1]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[2]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[3]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[4]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[5]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[6]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[7]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[8]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[9]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[10]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[11]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[12]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[13]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[14]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[15]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[16]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[17]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[18]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[19]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[20]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[21]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[22]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[23]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[24]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[25]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[26]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[27]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[28]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[29]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[30]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_0_t[31]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[0]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[1]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[2]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[3]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[4]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[5]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[6]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[7]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[8]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[9]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[10]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[11]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[12]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[13]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[14]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[15]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[16]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[17]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[18]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[19]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[20]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[21]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[22]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[23]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[24]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[25]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[26]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[27]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[28]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[29]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[30]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_1_t[31]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[0]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[1]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[2]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[3]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[4]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[5]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[6]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[7]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[8]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[9]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[10]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[11]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[12]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[13]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[14]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[15]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[16]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[17]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[18]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[19]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[20]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[21]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[22]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[23]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[24]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[25]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[26]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[27]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[28]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[29]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[30]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_4_t[31]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[0]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[1]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[2]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[3]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[4]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[5]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[6]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[7]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[8]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[9]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[10]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[11]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[12]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[13]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[14]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[15]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[16]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[17]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[18]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[19]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[20]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[21]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[22]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[23]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[24]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[25]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[26]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[27]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[28]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[29]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[30]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_5_t[31]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[0]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[1]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[2]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[3]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[4]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[5]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[6]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[7]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[8]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[9]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[10]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[11]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[12]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[13]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[14]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[15]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[16]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[17]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[18]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[19]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[20]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[21]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[22]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[23]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[24]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[25]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[26]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[27]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[28]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[29]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[30]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_6_t[31]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[0]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[1]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[2]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[3]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[4]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[5]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[6]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[7]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[8]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[9]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[10]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[11]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[12]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[13]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[14]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[15]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[16]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[17]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[18]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[19]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[20]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[21]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[22]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[23]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[24]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[25]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[26]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[27]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[28]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[29]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[30]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_7_t[31]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[0]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[1]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[2]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[3]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[4]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[5]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[6]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[7]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[8]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[9]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[10]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[11]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[12]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[13]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[14]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[15]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[16]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[17]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[18]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[19]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[20]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[21]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[22]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[23]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[24]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[25]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[26]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[27]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[28]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[29]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[30]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_8_t[31]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[0]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[1]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[2]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[3]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[4]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[5]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[6]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[7]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[8]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[9]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[10]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[11]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[12]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[13]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[14]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[15]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[16]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[17]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[18]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[19]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[20]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[21]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[22]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[23]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[24]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[25]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[26]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[27]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[28]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[29]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[30]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_15_t[31]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[0]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[1]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[2]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[3]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[4]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[5]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[6]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[7]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[8]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[9]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[10]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[11]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[12]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[13]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[14]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[15]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[16]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[17]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[18]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[19]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[20]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[21]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[22]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[23]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[24]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[25]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[26]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[27]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[28]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[29]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[30]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(regs_20_t[31]); // @[src/main/scala/device/AXI4DummySD.scala 72:43]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[0]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[1]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[2]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[3]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[4]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[5]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[6]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[7]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[8]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[9]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[10]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[11]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[12]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[13]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[14]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[15]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[16]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[17]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[18]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[19]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[20]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[21]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[22]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[23]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[24]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[25]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[26]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[27]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[28]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[29]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[30]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[31]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[32]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[33]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[34]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[35]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[36]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[37]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[38]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[39]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[40]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[41]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[42]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[43]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[44]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[45]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[46]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[47]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[48]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[49]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[50]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[51]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[52]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[53]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[54]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[55]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[56]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[57]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[58]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[59]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[60]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[61]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[62]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_REG_t[63]); // @[src/main/scala/device/AXI4DummySD.scala 144:44]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[0]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[1]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[2]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[3]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[4]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[5]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[6]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[7]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[8]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[9]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[10]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[11]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[12]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[13]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[14]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[15]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[16]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[17]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[18]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[19]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[20]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[21]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[22]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[23]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[24]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[25]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[26]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[27]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[28]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[29]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[30]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[31]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[32]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[33]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[34]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[35]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[36]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[37]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[38]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[39]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[40]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[41]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[42]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[43]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[44]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[45]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[46]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[47]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[48]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[49]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[50]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[51]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[52]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[53]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[54]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[55]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[56]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[57]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[58]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[59]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[60]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[61]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[62]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
    //
    if (enToggle_past) begin
      cover(io_in_r_bits_data_r_t[63]); // @[src/main/scala/device/AXI4DummySD.scala 144:36]
    end
  end
endmodule
module SimpleBus2AXI4Converter_3(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_resp_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_aw_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_out_w_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_w_bits_strb, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_b_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_ar_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_r_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_out_r_bits_data // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  toAXI4Lite = ~(io_in_req_valid & io_in_req_bits_cmd[1]); // @[src/main/scala/bus/simplebus/ToAXI4.scala 151:20]
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 | awAck & wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 189:53]
  wire  _GEN_2 = _wSend_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wen_T_1 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  _io_out_ar_valid_T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _io_out_aw_valid_T_1 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  wire  _io_out_w_valid_T_2 = ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:36]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  awAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  awAck_t = awAck ^ awAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_11668_clock;
  wire  toggle_11668_reset;
  wire  toggle_11668_valid;
  reg  toggle_11668_valid_reg;
  reg  wAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wAck_t = wAck ^ wAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_11669_clock;
  wire  toggle_11669_reset;
  wire  toggle_11669_valid;
  reg  toggle_11669_valid_reg;
  reg  wen_p; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  wen_t = wen ^ wen_p; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  toggle_11670_clock;
  wire  toggle_11670_reset;
  wire  toggle_11670_valid;
  reg  toggle_11670_valid_reg;
  GEN_w1_toggle #(.COVER_INDEX(11668)) toggle_11668 (
    .clock(toggle_11668_clock),
    .reset(toggle_11668_reset),
    .valid(toggle_11668_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(11669)) toggle_11669 (
    .clock(toggle_11669_clock),
    .reset(toggle_11669_reset),
    .valid(toggle_11669_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(11670)) toggle_11670 (
    .clock(toggle_11670_clock),
    .reset(toggle_11670_reset),
    .valid(toggle_11670_valid)
  );
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _io_out_w_valid_T_2 & io_out_w_ready : io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 199:25]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 183:23]
  assign io_out_aw_valid = _io_out_aw_valid_T_1 & ~awAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 193:33]
  assign io_out_aw_bits_addr = io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_w_valid = _io_out_aw_valid_T_1 & ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:33]
  assign io_out_w_bits_data = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 160:10]
  assign io_out_w_bits_strb = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 161:10]
  assign io_out_b_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 198:16]
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 158:12]
  assign io_out_r_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 197:16]
  assign toggle_11668_clock = clock;
  assign toggle_11668_reset = reset;
  assign toggle_11668_valid = awAck ^ toggle_11668_valid_reg;
  assign toggle_11669_clock = clock;
  assign toggle_11669_reset = reset;
  assign toggle_11669_valid = wAck ^ toggle_11669_valid_reg;
  assign toggle_11670_clock = clock;
  assign toggle_11670_reset = reset;
  assign toggle_11670_valid = wen ^ toggle_11670_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_2;
    end
    if (_wen_T_1) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
      wen <= io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~toAXI4Lite) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    awAck_p <= awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_11668_valid_reg <= awAck;
    wAck_p <= wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_11669_valid_reg <= wAck;
    wen_p <= wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    toggle_11670_valid_reg <= wen;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  awAck_p = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  toggle_11668_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  wAck_p = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  toggle_11669_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  wen_p = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  toggle_11670_valid_reg = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(toAXI4Lite); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
    end
    //
    if (enToggle_past) begin
      cover(awAck_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(wAck_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(wen_t); // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
  end
endmodule
module SimpleBus2AXI4Converter_4(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_resp_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_aw_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_out_w_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_w_bits_strb, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_b_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_r_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_valid // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  toAXI4Lite = ~(io_in_req_valid & io_in_req_bits_cmd[1]); // @[src/main/scala/bus/simplebus/ToAXI4.scala 151:20]
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 | awAck & wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 189:53]
  wire  _GEN_2 = _wSend_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wen_T_1 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  _io_out_ar_valid_T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _io_out_aw_valid_T_1 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  wire  _io_out_w_valid_T_2 = ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:36]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  awAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  awAck_t = awAck ^ awAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_11671_clock;
  wire  toggle_11671_reset;
  wire  toggle_11671_valid;
  reg  toggle_11671_valid_reg;
  reg  wAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wAck_t = wAck ^ wAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_11672_clock;
  wire  toggle_11672_reset;
  wire  toggle_11672_valid;
  reg  toggle_11672_valid_reg;
  reg  wen_p; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  wen_t = wen ^ wen_p; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  toggle_11673_clock;
  wire  toggle_11673_reset;
  wire  toggle_11673_valid;
  reg  toggle_11673_valid_reg;
  GEN_w1_toggle #(.COVER_INDEX(11671)) toggle_11671 (
    .clock(toggle_11671_clock),
    .reset(toggle_11671_reset),
    .valid(toggle_11671_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(11672)) toggle_11672 (
    .clock(toggle_11672_clock),
    .reset(toggle_11672_reset),
    .valid(toggle_11672_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(11673)) toggle_11673 (
    .clock(toggle_11673_clock),
    .reset(toggle_11673_reset),
    .valid(toggle_11673_valid)
  );
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _io_out_w_valid_T_2 & io_out_w_ready : 1'h1; // @[src/main/scala/bus/simplebus/ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 199:25]
  assign io_out_aw_valid = _io_out_aw_valid_T_1 & ~awAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 193:33]
  assign io_out_aw_bits_addr = io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_w_valid = _io_out_aw_valid_T_1 & ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:33]
  assign io_out_w_bits_data = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 160:10]
  assign io_out_w_bits_strb = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 161:10]
  assign io_out_b_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 198:16]
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 158:12]
  assign io_out_r_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 197:16]
  assign toggle_11671_clock = clock;
  assign toggle_11671_reset = reset;
  assign toggle_11671_valid = awAck ^ toggle_11671_valid_reg;
  assign toggle_11672_clock = clock;
  assign toggle_11672_reset = reset;
  assign toggle_11672_valid = wAck ^ toggle_11672_valid_reg;
  assign toggle_11673_clock = clock;
  assign toggle_11673_reset = reset;
  assign toggle_11673_valid = wen ^ toggle_11673_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_2;
    end
    if (_wen_T_1) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
      wen <= io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~toAXI4Lite) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    awAck_p <= awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_11671_valid_reg <= awAck;
    wAck_p <= wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_11672_valid_reg <= wAck;
    wen_p <= wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    toggle_11673_valid_reg <= wen;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  awAck_p = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  toggle_11671_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  wAck_p = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  toggle_11672_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  wen_p = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  toggle_11673_valid_reg = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(toAXI4Lite); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
    end
    //
    if (enToggle_past) begin
      cover(awAck_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(wAck_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(wen_t); // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
  end
endmodule
module SimpleBus2AXI4Converter_5(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_resp_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_b_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_ar_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_r_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_out_r_bits_data // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  toAXI4Lite = ~(io_in_req_valid & io_in_req_bits_cmd[1]); // @[src/main/scala/bus/simplebus/ToAXI4.scala 151:20]
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 | awAck & wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 189:53]
  wire  _GEN_2 = _wSend_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wen_T_1 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  _io_out_ar_valid_T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _io_out_aw_valid_T_1 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  wire  _io_out_w_valid_T_2 = ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:36]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  awAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  awAck_t = awAck ^ awAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_11674_clock;
  wire  toggle_11674_reset;
  wire  toggle_11674_valid;
  reg  toggle_11674_valid_reg;
  reg  wAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wAck_t = wAck ^ wAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_11675_clock;
  wire  toggle_11675_reset;
  wire  toggle_11675_valid;
  reg  toggle_11675_valid_reg;
  reg  wen_p; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  wen_t = wen ^ wen_p; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  toggle_11676_clock;
  wire  toggle_11676_reset;
  wire  toggle_11676_valid;
  reg  toggle_11676_valid_reg;
  GEN_w1_toggle #(.COVER_INDEX(11674)) toggle_11674 (
    .clock(toggle_11674_clock),
    .reset(toggle_11674_reset),
    .valid(toggle_11674_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(11675)) toggle_11675 (
    .clock(toggle_11675_clock),
    .reset(toggle_11675_reset),
    .valid(toggle_11675_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(11676)) toggle_11676 (
    .clock(toggle_11676_clock),
    .reset(toggle_11676_reset),
    .valid(toggle_11676_valid)
  );
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _io_out_w_valid_T_2 & io_out_w_ready : io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 199:25]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 183:23]
  assign io_out_aw_valid = _io_out_aw_valid_T_1 & ~awAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 193:33]
  assign io_out_w_valid = _io_out_aw_valid_T_1 & ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:33]
  assign io_out_b_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 198:16]
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 158:12]
  assign io_out_r_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 197:16]
  assign toggle_11674_clock = clock;
  assign toggle_11674_reset = reset;
  assign toggle_11674_valid = awAck ^ toggle_11674_valid_reg;
  assign toggle_11675_clock = clock;
  assign toggle_11675_reset = reset;
  assign toggle_11675_valid = wAck ^ toggle_11675_valid_reg;
  assign toggle_11676_clock = clock;
  assign toggle_11676_reset = reset;
  assign toggle_11676_valid = wen ^ toggle_11676_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_2;
    end
    if (_wen_T_1) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
      wen <= io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~toAXI4Lite) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    awAck_p <= awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_11674_valid_reg <= awAck;
    wAck_p <= wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_11675_valid_reg <= wAck;
    wen_p <= wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    toggle_11676_valid_reg <= wen;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  awAck_p = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  toggle_11674_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  wAck_p = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  toggle_11675_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  wen_p = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  toggle_11676_valid_reg = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(toAXI4Lite); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
    end
    //
    if (enToggle_past) begin
      cover(awAck_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(wAck_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(wen_t); // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
  end
endmodule
module SimpleBus2AXI4Converter_6(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_resp_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_b_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_ar_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_r_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_out_r_bits_data // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  toAXI4Lite = ~(io_in_req_valid & io_in_req_bits_cmd[1]); // @[src/main/scala/bus/simplebus/ToAXI4.scala 151:20]
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 | awAck & wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 189:53]
  wire  _GEN_2 = _wSend_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wen_T_1 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  _io_out_ar_valid_T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _io_out_aw_valid_T_1 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  wire  _io_out_w_valid_T_2 = ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:36]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  awAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  awAck_t = awAck ^ awAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_11677_clock;
  wire  toggle_11677_reset;
  wire  toggle_11677_valid;
  reg  toggle_11677_valid_reg;
  reg  wAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wAck_t = wAck ^ wAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_11678_clock;
  wire  toggle_11678_reset;
  wire  toggle_11678_valid;
  reg  toggle_11678_valid_reg;
  reg  wen_p; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  wen_t = wen ^ wen_p; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  toggle_11679_clock;
  wire  toggle_11679_reset;
  wire  toggle_11679_valid;
  reg  toggle_11679_valid_reg;
  GEN_w1_toggle #(.COVER_INDEX(11677)) toggle_11677 (
    .clock(toggle_11677_clock),
    .reset(toggle_11677_reset),
    .valid(toggle_11677_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(11678)) toggle_11678 (
    .clock(toggle_11678_clock),
    .reset(toggle_11678_reset),
    .valid(toggle_11678_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(11679)) toggle_11679 (
    .clock(toggle_11679_clock),
    .reset(toggle_11679_reset),
    .valid(toggle_11679_valid)
  );
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _io_out_w_valid_T_2 & io_out_w_ready : io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 199:25]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 183:23]
  assign io_out_aw_valid = _io_out_aw_valid_T_1 & ~awAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 193:33]
  assign io_out_w_valid = _io_out_aw_valid_T_1 & ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:33]
  assign io_out_b_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 198:16]
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 158:12]
  assign io_out_r_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 197:16]
  assign toggle_11677_clock = clock;
  assign toggle_11677_reset = reset;
  assign toggle_11677_valid = awAck ^ toggle_11677_valid_reg;
  assign toggle_11678_clock = clock;
  assign toggle_11678_reset = reset;
  assign toggle_11678_valid = wAck ^ toggle_11678_valid_reg;
  assign toggle_11679_clock = clock;
  assign toggle_11679_reset = reset;
  assign toggle_11679_valid = wen ^ toggle_11679_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_2;
    end
    if (_wen_T_1) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
      wen <= io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~toAXI4Lite) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    awAck_p <= awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_11677_valid_reg <= awAck;
    wAck_p <= wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_11678_valid_reg <= wAck;
    wen_p <= wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    toggle_11679_valid_reg <= wen;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  awAck_p = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  toggle_11677_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  wAck_p = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  toggle_11678_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  wen_p = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  toggle_11679_valid_reg = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(toAXI4Lite); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
    end
    //
    if (enToggle_past) begin
      cover(awAck_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(wAck_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(wen_t); // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
  end
endmodule
module SimpleBus2AXI4Converter_7(
  input         clock,
  input         reset,
  output        io_in_req_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_req_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [31:0] io_in_req_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [3:0]  io_in_req_bits_cmd, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [7:0]  io_in_req_bits_wmask, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_in_req_bits_wdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_in_resp_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_in_resp_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_in_resp_bits_rdata, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_aw_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_aw_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_aw_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_w_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_w_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [63:0] io_out_w_bits_data, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [7:0]  io_out_w_bits_strb, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_b_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_b_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_ar_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_ar_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output [31:0] io_out_ar_bits_addr, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  output        io_out_r_ready, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input         io_out_r_valid, // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
  input  [63:0] io_out_r_bits_data // @[src/main/scala/bus/simplebus/ToAXI4.scala 146:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  toAXI4Lite = ~(io_in_req_valid & io_in_req_bits_cmd[1]); // @[src/main/scala/bus/simplebus/ToAXI4.scala 151:20]
  wire  _awAck_T = io_out_aw_ready & io_out_aw_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  _GEN_0 = _awAck_T | awAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wSend_T_1 = io_out_w_ready & io_out_w_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wSend = _awAck_T & _wSend_T_1 | awAck & wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 189:53]
  wire  _GEN_2 = _wSend_T_1 | wAck; // @[src/main/scala/utils/StopWatch.scala 24:20 30:{20,24}]
  wire  _wen_T_1 = io_in_req_ready & io_in_req_valid; // @[src/main/scala/chisel3/util/Decoupled.scala 57:35]
  reg  wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  _io_out_ar_valid_T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 73:26]
  wire  _io_out_aw_valid_T_1 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/SimpleBus.scala 103:29]
  wire  _io_out_w_valid_T_2 = ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:36]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg  awAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  awAck_t = awAck ^ awAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_11680_clock;
  wire  toggle_11680_reset;
  wire  toggle_11680_valid;
  reg  toggle_11680_valid_reg;
  reg  wAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  wAck_t = wAck ^ wAck_p; // @[src/main/scala/utils/StopWatch.scala 24:20]
  wire  toggle_11681_clock;
  wire  toggle_11681_reset;
  wire  toggle_11681_valid;
  reg  toggle_11681_valid_reg;
  reg  wen_p; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  wen_t = wen ^ wen_p; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
  wire  toggle_11682_clock;
  wire  toggle_11682_reset;
  wire  toggle_11682_valid;
  reg  toggle_11682_valid_reg;
  GEN_w1_toggle #(.COVER_INDEX(11680)) toggle_11680 (
    .clock(toggle_11680_clock),
    .reset(toggle_11680_reset),
    .valid(toggle_11680_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(11681)) toggle_11681 (
    .clock(toggle_11681_clock),
    .reset(toggle_11681_reset),
    .valid(toggle_11681_valid)
  );
  GEN_w1_toggle #(.COVER_INDEX(11682)) toggle_11682 (
    .clock(toggle_11682_clock),
    .reset(toggle_11682_reset),
    .valid(toggle_11682_valid)
  );
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _io_out_w_valid_T_2 & io_out_w_ready : io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 199:25]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 183:23]
  assign io_out_aw_valid = _io_out_aw_valid_T_1 & ~awAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 193:33]
  assign io_out_aw_bits_addr = io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 182:6]
  assign io_out_w_valid = _io_out_aw_valid_T_1 & ~wAck; // @[src/main/scala/bus/simplebus/ToAXI4.scala 194:33]
  assign io_out_w_bits_data = io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 160:10]
  assign io_out_w_bits_strb = io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 161:10]
  assign io_out_b_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 198:16]
  assign io_out_ar_valid = io_in_req_valid & _io_out_ar_valid_T_4; // @[src/main/scala/bus/simplebus/SimpleBus.scala 104:29]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 158:12]
  assign io_out_r_ready = io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 197:16]
  assign toggle_11680_clock = clock;
  assign toggle_11680_reset = reset;
  assign toggle_11680_valid = awAck ^ toggle_11680_valid_reg;
  assign toggle_11681_clock = clock;
  assign toggle_11681_reset = reset;
  assign toggle_11681_valid = wAck ^ toggle_11681_valid_reg;
  assign toggle_11682_clock = clock;
  assign toggle_11682_reset = reset;
  assign toggle_11682_valid = wen ^ toggle_11682_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      awAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin // @[src/main/scala/utils/StopWatch.scala 24:20]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 24:20]
    end else if (wSend) begin // @[src/main/scala/utils/StopWatch.scala 31:19]
      wAck <= 1'h0; // @[src/main/scala/utils/StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_2;
    end
    if (_wen_T_1) begin // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
      wen <= io_in_req_bits_cmd[0]; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~toAXI4Lite) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    awAck_p <= awAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_11680_valid_reg <= awAck;
    wAck_p <= wAck; // @[src/main/scala/utils/StopWatch.scala 24:20]
    toggle_11681_valid_reg <= wAck;
    wen_p <= wen; // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    toggle_11682_valid_reg <= wen;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  awAck_p = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  toggle_11680_valid_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  wAck_p = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  toggle_11681_valid_reg = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  wen_p = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  toggle_11682_valid_reg = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(toAXI4Lite); // @[src/main/scala/bus/simplebus/ToAXI4.scala 153:9]
    end
    //
    if (enToggle_past) begin
      cover(awAck_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(wAck_t); // @[src/main/scala/utils/StopWatch.scala 24:20]
    end
    //
    if (enToggle_past) begin
      cover(wen_t); // @[src/main/scala/bus/simplebus/ToAXI4.scala 190:22]
    end
  end
endmodule
module SimMMIO(
  input         clock,
  input         reset,
  output        io_rw_req_ready, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input         io_rw_req_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [31:0] io_rw_req_bits_addr, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [3:0]  io_rw_req_bits_cmd, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [7:0]  io_rw_req_bits_wmask, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [63:0] io_rw_req_bits_wdata, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input         io_rw_resp_ready, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output        io_rw_resp_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output [3:0]  io_rw_resp_bits_cmd, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output [63:0] io_rw_resp_bits_rdata, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output        io_uart_out_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output [7:0]  io_uart_out_ch, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  output        io_uart_in_valid, // @[src/main/scala/sim/SimMMIO.scala 28:14]
  input  [7:0]  io_uart_in_ch // @[src/main/scala/sim/SimMMIO.scala 28:14]
);
  wire  xbar_clock; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_reset; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_in_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_in_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_in_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_in_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [7:0] xbar_io_in_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_in_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_in_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_in_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_in_resp_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_in_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_0_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_0_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_0_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_0_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_0_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_0_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_0_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_0_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_0_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_1_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_1_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_1_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_1_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_1_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_1_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_1_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_1_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_2_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_2_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_2_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_2_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_2_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_2_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_2_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_3_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_3_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_3_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_3_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_3_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_3_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_3_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_4_req_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_4_req_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_4_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_4_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_4_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_4_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_4_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  xbar_io_out_4_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_4_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 45:20]
  wire  uart_clock; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_reset; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [31:0] uart_io_in_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_w_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [63:0] uart_io_in_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [7:0] uart_io_in_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_b_ready; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [31:0] uart_io_in_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_r_ready; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [63:0] uart_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_extra_out_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [7:0] uart_io_extra_out_ch; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  uart_io_extra_in_valid; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire [7:0] uart_io_extra_in_ch; // @[src/main/scala/sim/SimMMIO.scala 48:20]
  wire  vga_clock; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_reset; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire [31:0] vga_io_in_fb_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_w_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_w_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire [63:0] vga_io_in_fb_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire [7:0] vga_io_in_fb_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_b_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_b_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_r_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_fb_r_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_w_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_w_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_b_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_b_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire [31:0] vga_io_in_ctrl_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_r_ready; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_r_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire [63:0] vga_io_in_ctrl_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  vga_io_vga_valid; // @[src/main/scala/sim/SimMMIO.scala 49:19]
  wire  flash_clock; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_reset; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_w_valid; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_b_ready; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire [31:0] flash_io_in_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_r_ready; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  flash_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire [63:0] flash_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 50:21]
  wire  sd_clock; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_reset; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire [31:0] sd_io_in_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_w_valid; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire [63:0] sd_io_in_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire [7:0] sd_io_in_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_b_ready; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire [31:0] sd_io_in_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_r_ready; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  sd_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire [63:0] sd_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 51:18]
  wire  uart_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] uart_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] uart_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] uart_io_in_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] uart_io_in_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] uart_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] uart_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] uart_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] uart_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] uart_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  uart_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] uart_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] vga_io_in_fb_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] vga_io_in_fb_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] vga_io_in_fb_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] vga_io_in_fb_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] vga_io_in_fb_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] vga_io_in_fb_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] vga_io_in_fb_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] vga_io_in_fb_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_fb_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] vga_io_in_ctrl_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] vga_io_in_ctrl_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] vga_io_in_ctrl_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] vga_io_in_ctrl_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  vga_io_in_ctrl_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] vga_io_in_ctrl_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] flash_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] flash_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] flash_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] flash_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  flash_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] flash_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_clock; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_reset; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_in_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] sd_io_in_bridge_io_in_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [3:0] sd_io_in_bridge_io_in_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] sd_io_in_bridge_io_in_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] sd_io_in_bridge_io_in_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_in_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] sd_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_aw_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_aw_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] sd_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_w_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_w_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] sd_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [7:0] sd_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_b_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_b_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_ar_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_ar_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [31:0] sd_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_r_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire  sd_io_in_bridge_io_out_r_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  wire [63:0] sd_io_in_bridge_io_out_r_bits_data; // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
  SimpleBusCrossbar1toN_1 xbar ( // @[src/main/scala/sim/SimMMIO.scala 45:20]
    .clock(xbar_clock),
    .reset(xbar_reset),
    .io_in_req_ready(xbar_io_in_req_ready),
    .io_in_req_valid(xbar_io_in_req_valid),
    .io_in_req_bits_addr(xbar_io_in_req_bits_addr),
    .io_in_req_bits_cmd(xbar_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(xbar_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(xbar_io_in_req_bits_wdata),
    .io_in_resp_ready(xbar_io_in_resp_ready),
    .io_in_resp_valid(xbar_io_in_resp_valid),
    .io_in_resp_bits_cmd(xbar_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(xbar_io_in_resp_bits_rdata),
    .io_out_0_req_ready(xbar_io_out_0_req_ready),
    .io_out_0_req_valid(xbar_io_out_0_req_valid),
    .io_out_0_req_bits_addr(xbar_io_out_0_req_bits_addr),
    .io_out_0_req_bits_cmd(xbar_io_out_0_req_bits_cmd),
    .io_out_0_req_bits_wmask(xbar_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wdata(xbar_io_out_0_req_bits_wdata),
    .io_out_0_resp_ready(xbar_io_out_0_resp_ready),
    .io_out_0_resp_valid(xbar_io_out_0_resp_valid),
    .io_out_0_resp_bits_rdata(xbar_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(xbar_io_out_1_req_ready),
    .io_out_1_req_valid(xbar_io_out_1_req_valid),
    .io_out_1_req_bits_addr(xbar_io_out_1_req_bits_addr),
    .io_out_1_req_bits_cmd(xbar_io_out_1_req_bits_cmd),
    .io_out_1_req_bits_wmask(xbar_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wdata(xbar_io_out_1_req_bits_wdata),
    .io_out_1_resp_ready(xbar_io_out_1_resp_ready),
    .io_out_1_resp_valid(xbar_io_out_1_resp_valid),
    .io_out_2_req_ready(xbar_io_out_2_req_ready),
    .io_out_2_req_valid(xbar_io_out_2_req_valid),
    .io_out_2_req_bits_addr(xbar_io_out_2_req_bits_addr),
    .io_out_2_req_bits_cmd(xbar_io_out_2_req_bits_cmd),
    .io_out_2_resp_ready(xbar_io_out_2_resp_ready),
    .io_out_2_resp_valid(xbar_io_out_2_resp_valid),
    .io_out_2_resp_bits_rdata(xbar_io_out_2_resp_bits_rdata),
    .io_out_3_req_ready(xbar_io_out_3_req_ready),
    .io_out_3_req_valid(xbar_io_out_3_req_valid),
    .io_out_3_req_bits_addr(xbar_io_out_3_req_bits_addr),
    .io_out_3_req_bits_cmd(xbar_io_out_3_req_bits_cmd),
    .io_out_3_resp_ready(xbar_io_out_3_resp_ready),
    .io_out_3_resp_valid(xbar_io_out_3_resp_valid),
    .io_out_3_resp_bits_rdata(xbar_io_out_3_resp_bits_rdata),
    .io_out_4_req_ready(xbar_io_out_4_req_ready),
    .io_out_4_req_valid(xbar_io_out_4_req_valid),
    .io_out_4_req_bits_addr(xbar_io_out_4_req_bits_addr),
    .io_out_4_req_bits_cmd(xbar_io_out_4_req_bits_cmd),
    .io_out_4_req_bits_wmask(xbar_io_out_4_req_bits_wmask),
    .io_out_4_req_bits_wdata(xbar_io_out_4_req_bits_wdata),
    .io_out_4_resp_ready(xbar_io_out_4_resp_ready),
    .io_out_4_resp_valid(xbar_io_out_4_resp_valid),
    .io_out_4_resp_bits_rdata(xbar_io_out_4_resp_bits_rdata)
  );
  AXI4UART uart ( // @[src/main/scala/sim/SimMMIO.scala 48:20]
    .clock(uart_clock),
    .reset(uart_reset),
    .io_in_aw_ready(uart_io_in_aw_ready),
    .io_in_aw_valid(uart_io_in_aw_valid),
    .io_in_aw_bits_addr(uart_io_in_aw_bits_addr),
    .io_in_w_ready(uart_io_in_w_ready),
    .io_in_w_valid(uart_io_in_w_valid),
    .io_in_w_bits_data(uart_io_in_w_bits_data),
    .io_in_w_bits_strb(uart_io_in_w_bits_strb),
    .io_in_b_ready(uart_io_in_b_ready),
    .io_in_b_valid(uart_io_in_b_valid),
    .io_in_ar_ready(uart_io_in_ar_ready),
    .io_in_ar_valid(uart_io_in_ar_valid),
    .io_in_ar_bits_addr(uart_io_in_ar_bits_addr),
    .io_in_r_ready(uart_io_in_r_ready),
    .io_in_r_valid(uart_io_in_r_valid),
    .io_in_r_bits_data(uart_io_in_r_bits_data),
    .io_extra_out_valid(uart_io_extra_out_valid),
    .io_extra_out_ch(uart_io_extra_out_ch),
    .io_extra_in_valid(uart_io_extra_in_valid),
    .io_extra_in_ch(uart_io_extra_in_ch)
  );
  AXI4VGA vga ( // @[src/main/scala/sim/SimMMIO.scala 49:19]
    .clock(vga_clock),
    .reset(vga_reset),
    .io_in_fb_aw_ready(vga_io_in_fb_aw_ready),
    .io_in_fb_aw_valid(vga_io_in_fb_aw_valid),
    .io_in_fb_aw_bits_addr(vga_io_in_fb_aw_bits_addr),
    .io_in_fb_w_ready(vga_io_in_fb_w_ready),
    .io_in_fb_w_valid(vga_io_in_fb_w_valid),
    .io_in_fb_w_bits_data(vga_io_in_fb_w_bits_data),
    .io_in_fb_w_bits_strb(vga_io_in_fb_w_bits_strb),
    .io_in_fb_b_ready(vga_io_in_fb_b_ready),
    .io_in_fb_b_valid(vga_io_in_fb_b_valid),
    .io_in_fb_ar_ready(vga_io_in_fb_ar_ready),
    .io_in_fb_ar_valid(vga_io_in_fb_ar_valid),
    .io_in_fb_r_ready(vga_io_in_fb_r_ready),
    .io_in_fb_r_valid(vga_io_in_fb_r_valid),
    .io_in_ctrl_aw_ready(vga_io_in_ctrl_aw_ready),
    .io_in_ctrl_aw_valid(vga_io_in_ctrl_aw_valid),
    .io_in_ctrl_w_ready(vga_io_in_ctrl_w_ready),
    .io_in_ctrl_w_valid(vga_io_in_ctrl_w_valid),
    .io_in_ctrl_b_ready(vga_io_in_ctrl_b_ready),
    .io_in_ctrl_b_valid(vga_io_in_ctrl_b_valid),
    .io_in_ctrl_ar_ready(vga_io_in_ctrl_ar_ready),
    .io_in_ctrl_ar_valid(vga_io_in_ctrl_ar_valid),
    .io_in_ctrl_ar_bits_addr(vga_io_in_ctrl_ar_bits_addr),
    .io_in_ctrl_r_ready(vga_io_in_ctrl_r_ready),
    .io_in_ctrl_r_valid(vga_io_in_ctrl_r_valid),
    .io_in_ctrl_r_bits_data(vga_io_in_ctrl_r_bits_data),
    .io_vga_valid(vga_io_vga_valid)
  );
  AXI4Flash flash ( // @[src/main/scala/sim/SimMMIO.scala 50:21]
    .clock(flash_clock),
    .reset(flash_reset),
    .io_in_aw_ready(flash_io_in_aw_ready),
    .io_in_aw_valid(flash_io_in_aw_valid),
    .io_in_w_ready(flash_io_in_w_ready),
    .io_in_w_valid(flash_io_in_w_valid),
    .io_in_b_ready(flash_io_in_b_ready),
    .io_in_b_valid(flash_io_in_b_valid),
    .io_in_ar_ready(flash_io_in_ar_ready),
    .io_in_ar_valid(flash_io_in_ar_valid),
    .io_in_ar_bits_addr(flash_io_in_ar_bits_addr),
    .io_in_r_ready(flash_io_in_r_ready),
    .io_in_r_valid(flash_io_in_r_valid),
    .io_in_r_bits_data(flash_io_in_r_bits_data)
  );
  AXI4DummySD sd ( // @[src/main/scala/sim/SimMMIO.scala 51:18]
    .clock(sd_clock),
    .reset(sd_reset),
    .io_in_aw_ready(sd_io_in_aw_ready),
    .io_in_aw_valid(sd_io_in_aw_valid),
    .io_in_aw_bits_addr(sd_io_in_aw_bits_addr),
    .io_in_w_ready(sd_io_in_w_ready),
    .io_in_w_valid(sd_io_in_w_valid),
    .io_in_w_bits_data(sd_io_in_w_bits_data),
    .io_in_w_bits_strb(sd_io_in_w_bits_strb),
    .io_in_b_ready(sd_io_in_b_ready),
    .io_in_b_valid(sd_io_in_b_valid),
    .io_in_ar_ready(sd_io_in_ar_ready),
    .io_in_ar_valid(sd_io_in_ar_valid),
    .io_in_ar_bits_addr(sd_io_in_ar_bits_addr),
    .io_in_r_ready(sd_io_in_r_ready),
    .io_in_r_valid(sd_io_in_r_valid),
    .io_in_r_bits_data(sd_io_in_r_bits_data)
  );
  SimpleBus2AXI4Converter_3 uart_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(uart_io_in_bridge_clock),
    .reset(uart_io_in_bridge_reset),
    .io_in_req_ready(uart_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(uart_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(uart_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(uart_io_in_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(uart_io_in_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(uart_io_in_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(uart_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(uart_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(uart_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(uart_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(uart_io_in_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(uart_io_in_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(uart_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(uart_io_in_bridge_io_out_w_valid),
    .io_out_w_bits_data(uart_io_in_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(uart_io_in_bridge_io_out_w_bits_strb),
    .io_out_b_ready(uart_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(uart_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(uart_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(uart_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(uart_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(uart_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(uart_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(uart_io_in_bridge_io_out_r_bits_data)
  );
  SimpleBus2AXI4Converter_4 vga_io_in_fb_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(vga_io_in_fb_bridge_clock),
    .reset(vga_io_in_fb_bridge_reset),
    .io_in_req_ready(vga_io_in_fb_bridge_io_in_req_ready),
    .io_in_req_valid(vga_io_in_fb_bridge_io_in_req_valid),
    .io_in_req_bits_addr(vga_io_in_fb_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(vga_io_in_fb_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(vga_io_in_fb_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(vga_io_in_fb_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(vga_io_in_fb_bridge_io_in_resp_ready),
    .io_in_resp_valid(vga_io_in_fb_bridge_io_in_resp_valid),
    .io_out_aw_ready(vga_io_in_fb_bridge_io_out_aw_ready),
    .io_out_aw_valid(vga_io_in_fb_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(vga_io_in_fb_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(vga_io_in_fb_bridge_io_out_w_ready),
    .io_out_w_valid(vga_io_in_fb_bridge_io_out_w_valid),
    .io_out_w_bits_data(vga_io_in_fb_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(vga_io_in_fb_bridge_io_out_w_bits_strb),
    .io_out_b_ready(vga_io_in_fb_bridge_io_out_b_ready),
    .io_out_b_valid(vga_io_in_fb_bridge_io_out_b_valid),
    .io_out_ar_valid(vga_io_in_fb_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(vga_io_in_fb_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(vga_io_in_fb_bridge_io_out_r_ready),
    .io_out_r_valid(vga_io_in_fb_bridge_io_out_r_valid)
  );
  SimpleBus2AXI4Converter_5 vga_io_in_ctrl_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(vga_io_in_ctrl_bridge_clock),
    .reset(vga_io_in_ctrl_bridge_reset),
    .io_in_req_ready(vga_io_in_ctrl_bridge_io_in_req_ready),
    .io_in_req_valid(vga_io_in_ctrl_bridge_io_in_req_valid),
    .io_in_req_bits_addr(vga_io_in_ctrl_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(vga_io_in_ctrl_bridge_io_in_req_bits_cmd),
    .io_in_resp_ready(vga_io_in_ctrl_bridge_io_in_resp_ready),
    .io_in_resp_valid(vga_io_in_ctrl_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(vga_io_in_ctrl_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(vga_io_in_ctrl_bridge_io_out_aw_ready),
    .io_out_aw_valid(vga_io_in_ctrl_bridge_io_out_aw_valid),
    .io_out_w_ready(vga_io_in_ctrl_bridge_io_out_w_ready),
    .io_out_w_valid(vga_io_in_ctrl_bridge_io_out_w_valid),
    .io_out_b_ready(vga_io_in_ctrl_bridge_io_out_b_ready),
    .io_out_b_valid(vga_io_in_ctrl_bridge_io_out_b_valid),
    .io_out_ar_ready(vga_io_in_ctrl_bridge_io_out_ar_ready),
    .io_out_ar_valid(vga_io_in_ctrl_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(vga_io_in_ctrl_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(vga_io_in_ctrl_bridge_io_out_r_ready),
    .io_out_r_valid(vga_io_in_ctrl_bridge_io_out_r_valid),
    .io_out_r_bits_data(vga_io_in_ctrl_bridge_io_out_r_bits_data)
  );
  SimpleBus2AXI4Converter_6 flash_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(flash_io_in_bridge_clock),
    .reset(flash_io_in_bridge_reset),
    .io_in_req_ready(flash_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(flash_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(flash_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(flash_io_in_bridge_io_in_req_bits_cmd),
    .io_in_resp_ready(flash_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(flash_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(flash_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(flash_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(flash_io_in_bridge_io_out_aw_valid),
    .io_out_w_ready(flash_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(flash_io_in_bridge_io_out_w_valid),
    .io_out_b_ready(flash_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(flash_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(flash_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(flash_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(flash_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(flash_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(flash_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(flash_io_in_bridge_io_out_r_bits_data)
  );
  SimpleBus2AXI4Converter_7 sd_io_in_bridge ( // @[src/main/scala/bus/simplebus/ToAXI4.scala 204:24]
    .clock(sd_io_in_bridge_clock),
    .reset(sd_io_in_bridge_reset),
    .io_in_req_ready(sd_io_in_bridge_io_in_req_ready),
    .io_in_req_valid(sd_io_in_bridge_io_in_req_valid),
    .io_in_req_bits_addr(sd_io_in_bridge_io_in_req_bits_addr),
    .io_in_req_bits_cmd(sd_io_in_bridge_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(sd_io_in_bridge_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(sd_io_in_bridge_io_in_req_bits_wdata),
    .io_in_resp_ready(sd_io_in_bridge_io_in_resp_ready),
    .io_in_resp_valid(sd_io_in_bridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(sd_io_in_bridge_io_in_resp_bits_rdata),
    .io_out_aw_ready(sd_io_in_bridge_io_out_aw_ready),
    .io_out_aw_valid(sd_io_in_bridge_io_out_aw_valid),
    .io_out_aw_bits_addr(sd_io_in_bridge_io_out_aw_bits_addr),
    .io_out_w_ready(sd_io_in_bridge_io_out_w_ready),
    .io_out_w_valid(sd_io_in_bridge_io_out_w_valid),
    .io_out_w_bits_data(sd_io_in_bridge_io_out_w_bits_data),
    .io_out_w_bits_strb(sd_io_in_bridge_io_out_w_bits_strb),
    .io_out_b_ready(sd_io_in_bridge_io_out_b_ready),
    .io_out_b_valid(sd_io_in_bridge_io_out_b_valid),
    .io_out_ar_ready(sd_io_in_bridge_io_out_ar_ready),
    .io_out_ar_valid(sd_io_in_bridge_io_out_ar_valid),
    .io_out_ar_bits_addr(sd_io_in_bridge_io_out_ar_bits_addr),
    .io_out_r_ready(sd_io_in_bridge_io_out_r_ready),
    .io_out_r_valid(sd_io_in_bridge_io_out_r_valid),
    .io_out_r_bits_data(sd_io_in_bridge_io_out_r_bits_data)
  );
  assign io_rw_req_ready = xbar_io_in_req_ready; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign io_rw_resp_valid = xbar_io_in_resp_valid; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign io_rw_resp_bits_cmd = xbar_io_in_resp_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign io_rw_resp_bits_rdata = xbar_io_in_resp_bits_rdata; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign io_uart_out_valid = uart_io_extra_out_valid; // @[src/main/scala/sim/SimMMIO.scala 65:21]
  assign io_uart_out_ch = uart_io_extra_out_ch; // @[src/main/scala/sim/SimMMIO.scala 65:21]
  assign io_uart_in_valid = uart_io_extra_in_valid; // @[src/main/scala/sim/SimMMIO.scala 65:21]
  assign xbar_clock = clock;
  assign xbar_reset = reset;
  assign xbar_io_in_req_valid = io_rw_req_valid; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_addr = io_rw_req_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_cmd = io_rw_req_bits_cmd; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_wmask = io_rw_req_bits_wmask; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_wdata = io_rw_req_bits_wdata; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_in_resp_ready = io_rw_resp_ready; // @[src/main/scala/sim/SimMMIO.scala 46:14]
  assign xbar_io_out_0_req_ready = uart_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_0_resp_valid = uart_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_0_resp_bits_rdata = uart_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_1_req_ready = vga_io_in_fb_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_1_resp_valid = vga_io_in_fb_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_2_req_ready = vga_io_in_ctrl_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_2_resp_valid = vga_io_in_ctrl_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_2_resp_bits_rdata = vga_io_in_ctrl_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_3_req_ready = flash_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_3_resp_valid = flash_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_3_resp_bits_rdata = flash_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_4_req_ready = sd_io_in_bridge_io_in_req_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_4_resp_valid = sd_io_in_bridge_io_in_resp_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign xbar_io_out_4_resp_bits_rdata = sd_io_in_bridge_io_in_resp_bits_rdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_clock = clock;
  assign uart_reset = reset;
  assign uart_io_in_aw_valid = uart_io_in_bridge_io_out_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_aw_bits_addr = uart_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_w_valid = uart_io_in_bridge_io_out_w_valid; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_w_bits_data = uart_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_w_bits_strb = uart_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_b_ready = uart_io_in_bridge_io_out_b_ready; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_ar_valid = uart_io_in_bridge_io_out_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_ar_bits_addr = uart_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_r_ready = uart_io_in_bridge_io_out_r_ready; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_extra_in_ch = io_uart_in_ch; // @[src/main/scala/sim/SimMMIO.scala 65:21]
  assign vga_clock = clock;
  assign vga_reset = reset;
  assign vga_io_in_fb_aw_valid = vga_io_in_fb_bridge_io_out_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_aw_bits_addr = vga_io_in_fb_bridge_io_out_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_w_valid = vga_io_in_fb_bridge_io_out_w_valid; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_w_bits_data = vga_io_in_fb_bridge_io_out_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_w_bits_strb = vga_io_in_fb_bridge_io_out_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_b_ready = vga_io_in_fb_bridge_io_out_b_ready; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_ar_valid = vga_io_in_fb_bridge_io_out_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_r_ready = vga_io_in_fb_bridge_io_out_r_ready; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_ctrl_aw_valid = vga_io_in_ctrl_bridge_io_out_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_w_valid = vga_io_in_ctrl_bridge_io_out_w_valid; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_b_ready = vga_io_in_ctrl_bridge_io_out_b_ready; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_ar_valid = vga_io_in_ctrl_bridge_io_out_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_ar_bits_addr = vga_io_in_ctrl_bridge_io_out_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_r_ready = vga_io_in_ctrl_bridge_io_out_r_ready; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign flash_clock = clock;
  assign flash_reset = reset;
  assign flash_io_in_aw_valid = flash_io_in_bridge_io_out_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_w_valid = flash_io_in_bridge_io_out_w_valid; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_b_ready = flash_io_in_bridge_io_out_b_ready; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_ar_valid = flash_io_in_bridge_io_out_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_ar_bits_addr = flash_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_r_ready = flash_io_in_bridge_io_out_r_ready; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign sd_clock = clock;
  assign sd_reset = reset;
  assign sd_io_in_aw_valid = sd_io_in_bridge_io_out_aw_valid; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_aw_bits_addr = sd_io_in_bridge_io_out_aw_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_w_valid = sd_io_in_bridge_io_out_w_valid; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_w_bits_data = sd_io_in_bridge_io_out_w_bits_data; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_w_bits_strb = sd_io_in_bridge_io_out_w_bits_strb; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_b_ready = sd_io_in_bridge_io_out_b_ready; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_ar_valid = sd_io_in_bridge_io_out_ar_valid; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_ar_bits_addr = sd_io_in_bridge_io_out_ar_bits_addr; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_r_ready = sd_io_in_bridge_io_out_r_ready; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign uart_io_in_bridge_clock = clock;
  assign uart_io_in_bridge_reset = reset;
  assign uart_io_in_bridge_io_in_req_valid = xbar_io_out_0_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_in_req_bits_addr = xbar_io_out_0_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_in_req_bits_cmd = xbar_io_out_0_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_in_req_bits_wmask = xbar_io_out_0_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_in_req_bits_wdata = xbar_io_out_0_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_in_resp_ready = xbar_io_out_0_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign uart_io_in_bridge_io_out_aw_ready = uart_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_bridge_io_out_w_ready = uart_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_bridge_io_out_b_valid = uart_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_bridge_io_out_ar_ready = uart_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_bridge_io_out_r_valid = uart_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign uart_io_in_bridge_io_out_r_bits_data = uart_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 54:14]
  assign vga_io_in_fb_bridge_clock = clock;
  assign vga_io_in_fb_bridge_reset = reset;
  assign vga_io_in_fb_bridge_io_in_req_valid = xbar_io_out_1_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_fb_bridge_io_in_req_bits_addr = xbar_io_out_1_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_fb_bridge_io_in_req_bits_cmd = xbar_io_out_1_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_fb_bridge_io_in_req_bits_wmask = xbar_io_out_1_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_fb_bridge_io_in_req_bits_wdata = xbar_io_out_1_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_fb_bridge_io_in_resp_ready = xbar_io_out_1_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_fb_bridge_io_out_aw_ready = vga_io_in_fb_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_bridge_io_out_w_ready = vga_io_in_fb_w_ready; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_bridge_io_out_b_valid = vga_io_in_fb_b_valid; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_fb_bridge_io_out_r_valid = vga_io_in_fb_r_valid; // @[src/main/scala/sim/SimMMIO.scala 55:16]
  assign vga_io_in_ctrl_bridge_clock = clock;
  assign vga_io_in_ctrl_bridge_reset = reset;
  assign vga_io_in_ctrl_bridge_io_in_req_valid = xbar_io_out_2_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_ctrl_bridge_io_in_req_bits_addr = xbar_io_out_2_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_ctrl_bridge_io_in_req_bits_cmd = xbar_io_out_2_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_ctrl_bridge_io_in_resp_ready = xbar_io_out_2_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign vga_io_in_ctrl_bridge_io_out_aw_ready = vga_io_in_ctrl_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_bridge_io_out_w_ready = vga_io_in_ctrl_w_ready; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_bridge_io_out_b_valid = vga_io_in_ctrl_b_valid; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_bridge_io_out_ar_ready = vga_io_in_ctrl_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_bridge_io_out_r_valid = vga_io_in_ctrl_r_valid; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign vga_io_in_ctrl_bridge_io_out_r_bits_data = vga_io_in_ctrl_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 56:18]
  assign flash_io_in_bridge_clock = clock;
  assign flash_io_in_bridge_reset = reset;
  assign flash_io_in_bridge_io_in_req_valid = xbar_io_out_3_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign flash_io_in_bridge_io_in_req_bits_addr = xbar_io_out_3_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign flash_io_in_bridge_io_in_req_bits_cmd = xbar_io_out_3_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign flash_io_in_bridge_io_in_resp_ready = xbar_io_out_3_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign flash_io_in_bridge_io_out_aw_ready = flash_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_bridge_io_out_w_ready = flash_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_bridge_io_out_b_valid = flash_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_bridge_io_out_ar_ready = flash_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_bridge_io_out_r_valid = flash_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign flash_io_in_bridge_io_out_r_bits_data = flash_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 57:15]
  assign sd_io_in_bridge_clock = clock;
  assign sd_io_in_bridge_reset = reset;
  assign sd_io_in_bridge_io_in_req_valid = xbar_io_out_4_req_valid; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign sd_io_in_bridge_io_in_req_bits_addr = xbar_io_out_4_req_bits_addr; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign sd_io_in_bridge_io_in_req_bits_cmd = xbar_io_out_4_req_bits_cmd; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign sd_io_in_bridge_io_in_req_bits_wmask = xbar_io_out_4_req_bits_wmask; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign sd_io_in_bridge_io_in_req_bits_wdata = xbar_io_out_4_req_bits_wdata; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign sd_io_in_bridge_io_in_resp_ready = xbar_io_out_4_resp_ready; // @[src/main/scala/bus/simplebus/ToAXI4.scala 205:18]
  assign sd_io_in_bridge_io_out_aw_ready = sd_io_in_aw_ready; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_bridge_io_out_w_ready = sd_io_in_w_ready; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_bridge_io_out_b_valid = sd_io_in_b_valid; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_bridge_io_out_ar_ready = sd_io_in_ar_ready; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_bridge_io_out_r_valid = sd_io_in_r_valid; // @[src/main/scala/sim/SimMMIO.scala 58:12]
  assign sd_io_in_bridge_io_out_r_bits_data = sd_io_in_r_bits_data; // @[src/main/scala/sim/SimMMIO.scala 58:12]
endmodule
module SimTop(
  input         reset,
  input         clock,
  output [63:0] difftest_exit, // @[difftest/src/main/scala/Difftest.scala 496:22]
  output [63:0] difftest_step, // @[difftest/src/main/scala/Difftest.scala 496:22]
  input         difftest_perfCtrl_clean, // @[difftest/src/main/scala/Difftest.scala 496:22]
  input         difftest_perfCtrl_dump, // @[difftest/src/main/scala/Difftest.scala 496:22]
  input  [63:0] difftest_logCtrl_begin, // @[difftest/src/main/scala/Difftest.scala 496:22]
  input  [63:0] difftest_logCtrl_end, // @[difftest/src/main/scala/Difftest.scala 496:22]
  input  [63:0] difftest_logCtrl_level, // @[difftest/src/main/scala/Difftest.scala 496:22]
  output        difftest_uart_out_valid, // @[difftest/src/main/scala/Difftest.scala 496:22]
  output [7:0]  difftest_uart_out_ch, // @[difftest/src/main/scala/Difftest.scala 496:22]
  output        difftest_uart_in_valid, // @[difftest/src/main/scala/Difftest.scala 496:22]
  input  [7:0]  difftest_uart_in_ch // @[difftest/src/main/scala/Difftest.scala 496:22]
);
assume property(reset == 1'b0);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  soc_clock; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_reset; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [31:0] soc_io_mem_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_w_ready; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_w_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [63:0] soc_io_mem_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [7:0] soc_io_mem_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_b_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [31:0] soc_io_mem_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [7:0] soc_io_mem_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [2:0] soc_io_mem_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_r_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [63:0] soc_io_mem_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mem_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mmio_req_ready; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mmio_req_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [31:0] soc_io_mmio_req_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [3:0] soc_io_mmio_req_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [7:0] soc_io_mmio_req_bits_wmask; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [63:0] soc_io_mmio_req_bits_wdata; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mmio_resp_ready; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  soc_io_mmio_resp_valid; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [3:0] soc_io_mmio_resp_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire [63:0] soc_io_mmio_resp_bits_rdata; // @[src/main/scala/sim/NutShellSim.scala 34:19]
  wire  mem_clock; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_reset; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [31:0] mem_io_in_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_w_ready; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_w_valid; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [63:0] mem_io_in_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [7:0] mem_io_in_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_b_valid; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_ar_ready; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [31:0] mem_io_in_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [7:0] mem_io_in_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [2:0] mem_io_in_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_r_valid; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire [63:0] mem_io_in_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  mem_io_in_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 35:19]
  wire  memdelay_clock; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_reset; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [31:0] memdelay_io_in_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_w_ready; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_w_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [63:0] memdelay_io_in_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [7:0] memdelay_io_in_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_b_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [31:0] memdelay_io_in_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [7:0] memdelay_io_in_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [2:0] memdelay_io_in_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_r_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [63:0] memdelay_io_in_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_in_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [31:0] memdelay_io_out_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_w_ready; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_w_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [63:0] memdelay_io_out_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [7:0] memdelay_io_out_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_b_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [31:0] memdelay_io_out_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [7:0] memdelay_io_out_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [2:0] memdelay_io_out_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_r_valid; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire [63:0] memdelay_io_out_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  memdelay_io_out_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 38:24]
  wire  mmio_clock; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_reset; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_io_rw_req_ready; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_io_rw_req_valid; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [31:0] mmio_io_rw_req_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [3:0] mmio_io_rw_req_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [7:0] mmio_io_rw_req_bits_wmask; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [63:0] mmio_io_rw_req_bits_wdata; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_io_rw_resp_ready; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_io_rw_resp_valid; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [3:0] mmio_io_rw_resp_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [63:0] mmio_io_rw_resp_bits_rdata; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_io_uart_out_valid; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [7:0] mmio_io_uart_out_ch; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire  mmio_io_uart_in_valid; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  wire [7:0] mmio_io_uart_in_ch; // @[src/main/scala/sim/NutShellSim.scala 39:20]
  reg [63:0] difftest_timer; // @[difftest/src/main/scala/Difftest.scala 501:24]
  wire [63:0] _difftest_timer_T_1 = difftest_timer + 64'h1; // @[difftest/src/main/scala/Difftest.scala 502:20]
  wire  difftest_log_enable = difftest_timer >= difftest_logCtrl_begin & difftest_timer < difftest_logCtrl_end; // @[difftest/src/main/scala/Difftest.scala 650:26]
  reg  enToggle = 1'h1;
  reg  enToggle_past = 1'h1;
  reg [63:0] difftest_timer_p; // @[difftest/src/main/scala/Difftest.scala 501:24]
  wire [63:0] difftest_timer_t = difftest_timer ^ difftest_timer_p; // @[difftest/src/main/scala/Difftest.scala 501:24]
  wire  toggle_11683_clock;
  wire  toggle_11683_reset;
  wire [63:0] toggle_11683_valid;
  reg [63:0] toggle_11683_valid_reg;
  NutShell soc ( // @[src/main/scala/sim/NutShellSim.scala 34:19]
    .clock(soc_clock),
    .reset(soc_reset),
    .io_mem_aw_ready(soc_io_mem_aw_ready),
    .io_mem_aw_valid(soc_io_mem_aw_valid),
    .io_mem_aw_bits_addr(soc_io_mem_aw_bits_addr),
    .io_mem_w_ready(soc_io_mem_w_ready),
    .io_mem_w_valid(soc_io_mem_w_valid),
    .io_mem_w_bits_data(soc_io_mem_w_bits_data),
    .io_mem_w_bits_strb(soc_io_mem_w_bits_strb),
    .io_mem_w_bits_last(soc_io_mem_w_bits_last),
    .io_mem_b_valid(soc_io_mem_b_valid),
    .io_mem_ar_valid(soc_io_mem_ar_valid),
    .io_mem_ar_bits_addr(soc_io_mem_ar_bits_addr),
    .io_mem_ar_bits_len(soc_io_mem_ar_bits_len),
    .io_mem_ar_bits_size(soc_io_mem_ar_bits_size),
    .io_mem_r_valid(soc_io_mem_r_valid),
    .io_mem_r_bits_data(soc_io_mem_r_bits_data),
    .io_mem_r_bits_last(soc_io_mem_r_bits_last),
    .io_mmio_req_ready(soc_io_mmio_req_ready),
    .io_mmio_req_valid(soc_io_mmio_req_valid),
    .io_mmio_req_bits_addr(soc_io_mmio_req_bits_addr),
    .io_mmio_req_bits_cmd(soc_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(soc_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(soc_io_mmio_req_bits_wdata),
    .io_mmio_resp_ready(soc_io_mmio_resp_ready),
    .io_mmio_resp_valid(soc_io_mmio_resp_valid),
    .io_mmio_resp_bits_cmd(soc_io_mmio_resp_bits_cmd),
    .io_mmio_resp_bits_rdata(soc_io_mmio_resp_bits_rdata)
  );
  AXI4RAM mem ( // @[src/main/scala/sim/NutShellSim.scala 35:19]
    .clock(mem_clock),
    .reset(mem_reset),
    .io_in_aw_ready(mem_io_in_aw_ready),
    .io_in_aw_valid(mem_io_in_aw_valid),
    .io_in_aw_bits_addr(mem_io_in_aw_bits_addr),
    .io_in_w_ready(mem_io_in_w_ready),
    .io_in_w_valid(mem_io_in_w_valid),
    .io_in_w_bits_data(mem_io_in_w_bits_data),
    .io_in_w_bits_strb(mem_io_in_w_bits_strb),
    .io_in_w_bits_last(mem_io_in_w_bits_last),
    .io_in_b_valid(mem_io_in_b_valid),
    .io_in_ar_ready(mem_io_in_ar_ready),
    .io_in_ar_valid(mem_io_in_ar_valid),
    .io_in_ar_bits_addr(mem_io_in_ar_bits_addr),
    .io_in_ar_bits_len(mem_io_in_ar_bits_len),
    .io_in_ar_bits_size(mem_io_in_ar_bits_size),
    .io_in_r_valid(mem_io_in_r_valid),
    .io_in_r_bits_data(mem_io_in_r_bits_data),
    .io_in_r_bits_last(mem_io_in_r_bits_last)
  );
  AXI4Delayer memdelay ( // @[src/main/scala/sim/NutShellSim.scala 38:24]
    .clock(memdelay_clock),
    .reset(memdelay_reset),
    .io_in_aw_ready(memdelay_io_in_aw_ready),
    .io_in_aw_valid(memdelay_io_in_aw_valid),
    .io_in_aw_bits_addr(memdelay_io_in_aw_bits_addr),
    .io_in_w_ready(memdelay_io_in_w_ready),
    .io_in_w_valid(memdelay_io_in_w_valid),
    .io_in_w_bits_data(memdelay_io_in_w_bits_data),
    .io_in_w_bits_strb(memdelay_io_in_w_bits_strb),
    .io_in_w_bits_last(memdelay_io_in_w_bits_last),
    .io_in_b_valid(memdelay_io_in_b_valid),
    .io_in_ar_valid(memdelay_io_in_ar_valid),
    .io_in_ar_bits_addr(memdelay_io_in_ar_bits_addr),
    .io_in_ar_bits_len(memdelay_io_in_ar_bits_len),
    .io_in_ar_bits_size(memdelay_io_in_ar_bits_size),
    .io_in_r_valid(memdelay_io_in_r_valid),
    .io_in_r_bits_data(memdelay_io_in_r_bits_data),
    .io_in_r_bits_last(memdelay_io_in_r_bits_last),
    .io_out_aw_ready(memdelay_io_out_aw_ready),
    .io_out_aw_valid(memdelay_io_out_aw_valid),
    .io_out_aw_bits_addr(memdelay_io_out_aw_bits_addr),
    .io_out_w_ready(memdelay_io_out_w_ready),
    .io_out_w_valid(memdelay_io_out_w_valid),
    .io_out_w_bits_data(memdelay_io_out_w_bits_data),
    .io_out_w_bits_strb(memdelay_io_out_w_bits_strb),
    .io_out_w_bits_last(memdelay_io_out_w_bits_last),
    .io_out_b_valid(memdelay_io_out_b_valid),
    .io_out_ar_valid(memdelay_io_out_ar_valid),
    .io_out_ar_bits_addr(memdelay_io_out_ar_bits_addr),
    .io_out_ar_bits_len(memdelay_io_out_ar_bits_len),
    .io_out_ar_bits_size(memdelay_io_out_ar_bits_size),
    .io_out_r_valid(memdelay_io_out_r_valid),
    .io_out_r_bits_data(memdelay_io_out_r_bits_data),
    .io_out_r_bits_last(memdelay_io_out_r_bits_last)
  );
  SimMMIO mmio ( // @[src/main/scala/sim/NutShellSim.scala 39:20]
    .clock(mmio_clock),
    .reset(mmio_reset),
    .io_rw_req_ready(mmio_io_rw_req_ready),
    .io_rw_req_valid(mmio_io_rw_req_valid),
    .io_rw_req_bits_addr(mmio_io_rw_req_bits_addr),
    .io_rw_req_bits_cmd(mmio_io_rw_req_bits_cmd),
    .io_rw_req_bits_wmask(mmio_io_rw_req_bits_wmask),
    .io_rw_req_bits_wdata(mmio_io_rw_req_bits_wdata),
    .io_rw_resp_ready(mmio_io_rw_resp_ready),
    .io_rw_resp_valid(mmio_io_rw_resp_valid),
    .io_rw_resp_bits_cmd(mmio_io_rw_resp_bits_cmd),
    .io_rw_resp_bits_rdata(mmio_io_rw_resp_bits_rdata),
    .io_uart_out_valid(mmio_io_uart_out_valid),
    .io_uart_out_ch(mmio_io_uart_out_ch),
    .io_uart_in_valid(mmio_io_uart_in_valid),
    .io_uart_in_ch(mmio_io_uart_in_ch)
  );
  GEN_w64_toggle #(.COVER_INDEX(11683)) toggle_11683 (
    .clock(toggle_11683_clock),
    .reset(toggle_11683_reset),
    .valid(toggle_11683_valid)
  );
  assign difftest_exit = 64'h0; // @[difftest/src/main/scala/Difftest.scala 498:19]
  assign difftest_step = 64'h1; // @[difftest/src/main/scala/Difftest.scala 499:19]
  assign difftest_uart_out_valid = mmio_io_uart_out_valid; // @[src/main/scala/sim/NutShellSim.scala 64:17]
  assign difftest_uart_out_ch = mmio_io_uart_out_ch; // @[src/main/scala/sim/NutShellSim.scala 64:17]
  assign difftest_uart_in_valid = mmio_io_uart_in_valid; // @[src/main/scala/sim/NutShellSim.scala 64:17]
  assign soc_clock = clock;
  assign soc_reset = reset;
  assign soc_io_mem_aw_ready = memdelay_io_in_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign soc_io_mem_w_ready = memdelay_io_in_w_ready; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign soc_io_mem_b_valid = memdelay_io_in_b_valid; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign soc_io_mem_r_valid = memdelay_io_in_r_valid; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign soc_io_mem_r_bits_data = memdelay_io_in_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign soc_io_mem_r_bits_last = memdelay_io_in_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign soc_io_mmio_req_ready = mmio_io_rw_req_ready; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign soc_io_mmio_resp_valid = mmio_io_rw_resp_valid; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign soc_io_mmio_resp_bits_cmd = mmio_io_rw_resp_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign soc_io_mmio_resp_bits_rdata = mmio_io_rw_resp_bits_rdata; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_io_in_aw_valid = memdelay_io_out_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_aw_bits_addr = memdelay_io_out_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_w_valid = memdelay_io_out_w_valid; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_w_bits_data = memdelay_io_out_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_w_bits_strb = memdelay_io_out_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_w_bits_last = memdelay_io_out_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_ar_valid = memdelay_io_out_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_ar_bits_addr = memdelay_io_out_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_ar_bits_len = memdelay_io_out_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mem_io_in_ar_bits_size = memdelay_io_out_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign memdelay_clock = clock;
  assign memdelay_reset = reset;
  assign memdelay_io_in_aw_valid = soc_io_mem_aw_valid; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_aw_bits_addr = soc_io_mem_aw_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_w_valid = soc_io_mem_w_valid; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_w_bits_data = soc_io_mem_w_bits_data; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_w_bits_strb = soc_io_mem_w_bits_strb; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_w_bits_last = soc_io_mem_w_bits_last; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_ar_valid = soc_io_mem_ar_valid; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_ar_bits_addr = soc_io_mem_ar_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_ar_bits_len = soc_io_mem_ar_bits_len; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_in_ar_bits_size = soc_io_mem_ar_bits_size; // @[src/main/scala/sim/NutShellSim.scala 43:18]
  assign memdelay_io_out_aw_ready = mem_io_in_aw_ready; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign memdelay_io_out_w_ready = mem_io_in_w_ready; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign memdelay_io_out_b_valid = mem_io_in_b_valid; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign memdelay_io_out_r_valid = mem_io_in_r_valid; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign memdelay_io_out_r_bits_data = mem_io_in_r_bits_data; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign memdelay_io_out_r_bits_last = mem_io_in_r_bits_last; // @[src/main/scala/sim/NutShellSim.scala 44:13]
  assign mmio_clock = clock;
  assign mmio_reset = reset;
  assign mmio_io_rw_req_valid = soc_io_mmio_req_valid; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mmio_io_rw_req_bits_addr = soc_io_mmio_req_bits_addr; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mmio_io_rw_req_bits_cmd = soc_io_mmio_req_bits_cmd; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mmio_io_rw_req_bits_wmask = soc_io_mmio_req_bits_wmask; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mmio_io_rw_req_bits_wdata = soc_io_mmio_req_bits_wdata; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mmio_io_rw_resp_ready = soc_io_mmio_resp_ready; // @[src/main/scala/sim/NutShellSim.scala 46:14]
  assign mmio_io_uart_in_ch = difftest_uart_in_ch; // @[src/main/scala/sim/NutShellSim.scala 64:17]
  assign toggle_11683_clock = clock;
  assign toggle_11683_reset = reset;
  assign toggle_11683_valid = difftest_timer ^ toggle_11683_valid_reg;
  always @(posedge clock) begin
    if (reset) begin // @[difftest/src/main/scala/Difftest.scala 501:24]
      difftest_timer <= 64'h0; // @[difftest/src/main/scala/Difftest.scala 501:24]
    end else begin
      difftest_timer <= _difftest_timer_T_1; // @[difftest/src/main/scala/Difftest.scala 502:11]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(difftest_logCtrl_begin <= difftest_logCtrl_end)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at NutShellSim.scala:57 assert(log_begin <= log_end)\n"); // @[src/main/scala/sim/NutShellSim.scala 57:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    enToggle <= 1'h1;
    enToggle_past <= enToggle;
    difftest_timer_p <= difftest_timer; // @[difftest/src/main/scala/Difftest.scala 501:24]
    toggle_11683_valid_reg <= difftest_timer;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  difftest_timer = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  difftest_timer_p = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  toggle_11683_valid_reg = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(difftest_logCtrl_begin <= difftest_logCtrl_end); // @[src/main/scala/sim/NutShellSim.scala 57:9]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[0]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[1]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[2]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[3]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[4]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[5]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[6]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[7]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[8]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[9]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[10]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[11]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[12]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[13]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[14]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[15]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[16]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[17]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[18]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[19]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[20]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[21]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[22]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[23]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[24]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[25]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[26]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[27]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[28]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[29]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[30]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[31]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[32]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[33]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[34]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[35]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[36]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[37]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[38]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[39]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[40]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[41]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[42]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[43]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[44]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[45]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[46]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[47]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[48]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[49]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[50]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[51]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[52]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[53]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[54]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[55]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[56]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[57]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[58]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[59]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[60]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[61]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[62]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
    //
    if (enToggle_past) begin
      cover(difftest_timer_t[63]); // @[difftest/src/main/scala/Difftest.scala 501:24]
    end
  end
endmodule
module array_0(
  input  [8:0]  R0_addr,
  input         R0_en,
  input         R0_clk,
  output [73:0] R0_data,
  input  [8:0]  W0_addr,
  input         W0_en,
  input         W0_clk,
  input  [73:0] W0_data
);
  wire [8:0] array_0_ext_R0_addr;
  wire  array_0_ext_R0_en;
  wire  array_0_ext_R0_clk;
  wire [73:0] array_0_ext_R0_data;
  wire [8:0] array_0_ext_W0_addr;
  wire  array_0_ext_W0_en;
  wire  array_0_ext_W0_clk;
  wire [73:0] array_0_ext_W0_data;
  array_0_ext array_0_ext (
    .R0_addr(array_0_ext_R0_addr),
    .R0_en(array_0_ext_R0_en),
    .R0_clk(array_0_ext_R0_clk),
    .R0_data(array_0_ext_R0_data),
    .W0_addr(array_0_ext_W0_addr),
    .W0_en(array_0_ext_W0_en),
    .W0_clk(array_0_ext_W0_clk),
    .W0_data(array_0_ext_W0_data)
  );
  assign array_0_ext_R0_clk = R0_clk;
  assign array_0_ext_R0_en = R0_en;
  assign array_0_ext_R0_addr = R0_addr;
  assign R0_data = array_0_ext_R0_data[73:0];
  assign array_0_ext_W0_clk = W0_clk;
  assign array_0_ext_W0_en = W0_en;
  assign array_0_ext_W0_addr = W0_addr;
  assign array_0_ext_W0_data = W0_data;
endmodule
